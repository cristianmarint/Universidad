��  CCircuit��  CSerializeHack           ��  CPart  H � H �     ���  CEarth�� 	 CTerminal  p�q�      @ 	         @A�c=�?    c�{�         ��      �� 
 CResistors��  CValue  Y �y �    220          �k@      �?   
�  � �� �      � 	 {��.@�W�/�1�?  
�  � �� �      � 	 {��.@�W�/�1�?  
�  � �� �      � 	 {��.@�W�/�1�?  
�  � �� �      � 	        �          
�  � �� �      � 	 {��.@�W�/�1�?  
�  � �� �      � 	 {��.@�W�/�1�?  
�  � �� �      � 	 {��.@�W�/�1�?  
�  � �� �      �          �          
�  � �� �     �          �          
�  � �� �     }   �i�n� @�W�/�1��  
�  � �� �     �   �i�n� @�W�/�1��  
�  � �� �     |   �i�n� @�W�/�1��  
�  � �� �     �          �          
�  � �� �     �   �i�n� @�W�/�1��  
�  � �� �     �   �i�n� @�W�/�1��  
�  � �� �     �   �i�n� @�W�/�1��    z �� �          �� v   ��  CSevenSegmentDisplay
�  � 0� 1     �          �          
�  � @� A     |   �i�n� @ W�/�1�?  
�  � P� Q     �   �i�n� @ W�/�1�?  
�  � `� a     }   �i�n� @ W�/�1�?  
�  � l� �     �           @A�c=岿  
�  � `� a     �          �          
�  � P� Q     �   �i�n� @ W�/�1�?  
�  � @� A     �   �i�n� @ W�/�1�?  
�  � 0� 1     �   �i�n� @ W�/�1�?    � ,� l     " 	     ��0 <           �
�  � �� �      � 	         @A�c=�?    � �� �     ,    ��       �
�  H8]9     D          �          
�  HH]I     E   �i�n� @ W�/�1�?  
�  HX]Y     F   �i�n� @ W�/�1�?  
�  Hh]i     G   �i�n� @ W�/�1�?  
�  ptq�     @           @A�c=岿  
�  �h�i     ?          �          
�  �X�Y     A   �i�n� @ W�/�1�?  
�  �H�I     B   �i�n� @ W�/�1�?  
�  �8�9     C   �i�n� @ W�/�1�?    \4�t     . 	     ��0 <           ��  	�)�    220          �k@      �?   
�  ����      J 	 {��.@�W�/�1�?  
�  ����      K 	 {��.@�W�/�1�?  
�  ����      L 	 {��.@�W�/�1�?  
�  p�q�      � 	        �          
�  `�a�      , 	 |��.@�W�/�1�?  
�  P�Q�      � 	 {��.@�W�/�1�?  
�  @�A�      � 	 {��.@�W�/�1�?  
�  0�1�      I          �          
�  0�1�     H          �          
�  @�A�     G   �i�n� @�W�/�1��  
�  P�Q�     F   �i�n� @�W�/�1��  
�  `�a�     E   �i�n� @�W�/�1��  
�  p�q�     D          �          
�  ����     C   �i�n� @�W�/�1��  
�  ����     B   �i�n� @�W�/�1��  
�  ����     A   �i�n� @�W�/�1��    *���    9      �� v   ��  C4511
�  �p��      �          �          
�  �p��      �          �          
�  �p��      �          �          
�  ppq�      �          �          
�  `pa�      �         @          
�  PpQ�      �         @          
�  @pA�      �          �          
�  @�A�     �   {��.@�W�/�1��  
�  P�Q�     �   {��.@�W�/�1��  
�  `�a�     ,   |��.@�W�/�1��  
�  p�q�     �          �          
�  ����     L   {��.@�W�/�1��  
�  ����     K   {��.@�W�/�1��  
�  ����     J   {��.@�W�/�1��    8���    K      ��  h   I�
�  � h� }      �          �          
�  � h� }      �          �          
�  � h� }      �          �          
�  � h� }      �          �          
�  � h� }      �         @          
�  � h� }      �         @          
�  � h� }      �          �          
�  � �� �     �   {��.@�W�/�1��  
�  � �� �     �   {��.@�W�/�1��  
�  � �� �     �   {��.@�W�/�1��  
�  � �� �     �          �          
�  � �� �     �   {��.@�W�/�1��  
�  � �� �     �   {��.@�W�/�1��  
�  � �� �     �   {��.@�W�/�1��    � |� �    Z      ��  h   �� 
 CCounter10
�  � �       �         @          
�  � �       �          �          
�  � 0� 1     �          �          
�  � <� Q     �          �          
�  � <� Q     �          �          
�  � <� Q     �          �          
�  � <� Q     �          �            � � <    j      ��  ,   h�
�  ��      �         @          
�  xy      �          �          
�  X0m1     �          �          
�  p<qQ     �          �          
�  �<�Q     �          �          
�  �<�Q     �          �          
�  �<�Q     �          �            l�<    r      ��  ,   ��  CAND
�  4HII     �          �          
�  48I9     �          �          
�  @A     �          �            44L    {      ��    y�
�  �H�I     �          �          
�  �8�9     �          �          
�  `@uA     �          �            t4�L          ��    h�
�  ��      �         @          
�  ��      ~          �          
�  �0�1     �          �          
�  �<�Q     �          �          
�  �<�Q     �          �          
�  �<�Q     �          �          
�  �<�Q     �          �            ��<    �      ��  ,   h�
�  @A      �         @          
�   !      �          �          
�   01     �          �          
�  <Q     �          �          
�  (<)Q     �          �          
�  8<9Q     �         @          
�  H<IQ     �          �            L<    �      ��  ,   I�
�  HhI}      �          �          
�  8h9}      �         @          
�  (h)}      �          �          
�  h}      �          �          
�  h	}      �         @          
�  �h�}      �         @          
�  �h�}      �          �          
�  ����     �   |��.@�W�/�1��  
�  ����     �   |��.@�W�/�1��  
�  �	�     �          �          
�  ��     �   |��.@�W�/�1��  
�  (�)�     �   |��.@�W�/�1��  
�  8�9�     �   |��.@�W�/�1��  
�  H�I�     �          �            �|L�    �      ��  h   I�
�  �p��      �          �          
�  �p��      �          �          
�  �p��      �          �          
�  �p��      �          �          
�  �p��      �         @          
�  �p��      �         @          
�  �p��      �          �          
�  ����     �   {��.@�W�/�1��  
�  ����     �   {��.@�W�/�1��  
�  ����     �   {��.@�W�/�1��  
�  ����     �          �          
�  ����     �   {��.@�W�/�1��  
�  ����     �   {��.@�W�/�1��  
�  ����     �   {��.@�W�/�1��    ����    �      ��  h   ��  a���    220          �k@      �?   
�  ����      � 	 {��.@�W�/�1�?  
�  ����      � 	 {��.@�W�/�1�?  
�  ����      � 	 {��.@�W�/�1�?  
�  ����      � 	        �          
�  ����      � 	 {��.@�W�/�1�?  
�  ����      � 	 {��.@�W�/�1�?  
�  ����      � 	 {��.@�W�/�1�?  
�  ����      �          �          
�  ����     �          �          
�  ����     �   �i�n� @�W�/�1��  
�  ����     �   �i�n� @�W�/�1��  
�  ����     �   �i�n� @�W�/�1��  
�  ����     �          �          
�  ����     �   �i�n� @�W�/�1��  
�  ����     �   �i�n� @�W�/�1��  
�  ����     �   �i�n� @�W�/�1��    ����    �      �� v    �
�  �8�9     �          �          
�  �H�I     �   �i�n� @ W�/�1�?  
�  �X�Y     �   �i�n� @ W�/�1�?  
�  �h�i     �   �i�n� @ W�/�1�?  
�  �t��     �           @A�c=岿  
�  �h�i     �          �          
�  �X�Y     �   �i�n� @ W�/�1�?  
�  �H�I     �   �i�n� @ W�/�1�?  
�  �8�9     �   �i�n� @ W�/�1�?    �4�t     � 	     ��0 <           �
�  ��      � 	         �l��~�?    �#�     �    ��       �
�  �01     �   �i�n� @ W�/�1�?  
�  �@A     �          �          
�  �PQ     �   �i�n� @ W�/�1�?  
�  �`a     �   �i�n� @ W�/�1�?  
�  l�     �           �l��~��  
�  4`Ia     �          �          
�  4PIQ     �          �          
�  4@IA     �   �i�n� @ W�/�1�?  
�  40I1     �   �i�n� @ W�/�1�?    ,4l     � 	     ��0 <             ��  ����    220          �k@      �?   
�  H�I�      � 	        �          
�  8�9�      � 	 |��.@�W�/�1�?  
�  (�)�      � 	 |��.@�W�/�1�?  
�  ��      � 	 |��.@�W�/�1�?  
�  �	�      � 	        �          
�  ����      � 	 |��.@�W�/�1�?  
�  ����      � 	 |��.@�W�/�1�?  
�  ����      �          �          
�  ����     �          �          
�  ����     �   �i�n� @�W�/�1��  
�  ����     �   �i�n� @�W�/�1��  
�  �	�     �          �          
�  ��     �   �i�n� @�W�/�1��  
�  (�)�     �   �i�n� @�W�/�1��  
�  8�9�     �   �i�n� @�W�/�1��  
�  H�I�     �          �            ��L�    �      �� v   �
�  ����      � 	         @A�c=�?    ����     �    ��      y�
�  �4�I     �         @          
�  �4�I     �          �          
�  ��      �          �            ��4    �      ��    y�
�  8$99     W          �          
�  H$I9               �          
�  @�A      ~          �            4L$    �      ��    ��  CBattery�  DGlU    5V         @      �? V 
�  d`ya     N         @          
�  8`Ma     O                       LTdl    �    ��      ��  CSPST��  CToggle  �h��     �   
�  x`�a     N 	       @          
�  �`�a     �         @            �\�d     �     ��    �
�  (x)�      ) 	         �l��~�?    �3�         ��      y�
�  � �      R         @          
�  � �      U         @          
�  �,�A     +         @            ��,         ��    ��  �1�    220          �k@      �?   
�  ����      _ 	 |��.@�W�/�1�?  
�  ����      ^ 	 |��.@�W�/�1�?  
�  ����      ] 	        �          
�  x�y�      \ 	        �          
�  h�i�      [ 	        �          
�  X�Y�      Z 	        �          
�  H�I�      Y 	        �          
�  8�9�      {          �          
�  8�9�     p          �          
�  H�I�     v          �          
�  X�Y�     u          �          
�  h�i�     t          �          
�  x�y�     s          �          
�  ����     z          �          
�  ����     y   �i�n� @�W�/�1��  
�  ����     x   �i�n� @�W�/�1��    2���         �� v    �
�  P e!     s          �          
�  P0e1     t          �          
�  P@eA     u          �          
�  PPeQ     v          �          
�  x\yq     r            W�/�1��  
�  �P�Q     w          �          
�  �@�A     x   �i�n� @ W�/�1�?  
�  �0�1     y   �i�n� @ W�/�1�?  
�  � �!     z          �            d�\     	     ��0 <             �
�  xpy�      r 	          W�/�1�?    k���     "   ��      �
�  ����     M            �:�?    �|�    $   ��       �
�   ()     l   �i�n� @ W�/�1�?  
�   89     k   �i�n� @ W�/�1�?  
�   HI     j          �          
�   XY     i          �          
�  (d)y     )           �l��~��  
�  DXYY     q          �          
�  DHYI     o   �i�n� @ W�/�1�?  
�  D8Y9     n   �i�n� @ W�/�1�?  
�  D(Y)     m   �i�n� @ W�/�1�?    $Dd     &	     ��0 <            ��  ����    220          �k@      �?   
�  X�Y�      f 	 |��.@�W�/�1�?  
�  H�I�      e 	 |��.@�W�/�1�?  
�  8�9�      d 	 |��.@�W�/�1�?  
�  (�)�      c 	 |��.@�W�/�1�?  
�  ��      b 	 |��.@�W�/�1�?  
�  �	�      a 	        �          
�  ����      ` 	        �          
�  ����      g          �          
�  ����     h          �          
�  ����     i          �          
�  �	�     j          �          
�  ��     k   �i�n� @�W�/�1��  
�  (�)�     l   �i�n� @�W�/�1��  
�  8�9�     m   �i�n� @�W�/�1��  
�  H�I�     n   �i�n� @�W�/�1��  
�  X�Y�     o   �i�n� @�W�/�1��    ��\�    1     �� v   I�
�  X`Yu      U         @          
�  H`Iu      T          �          
�  8`9u      S          �          
�  (`)u      R         @          
�  `u      �         @          
�  `	u      �         @          
�  �`�u      M                     
�  ����     `          �          
�  �	�     a          �          
�  ��     b   |��.@�W�/�1��  
�  (�)�     c   |��.@�W�/�1��  
�  8�9�     d   |��.@�W�/�1��  
�  H�I�     e   |��.@�W�/�1��  
�  X�Y�     f   |��.@�W�/�1��    �t\�    B     ��  h   I�
�  �X�m      X         @          
�  �X�m      W          �          
�  �X�m                �          
�  xXym      �          �          
�  hXim      �         @          
�  XXYm      �         @          
�  HXIm      M                     
�  H�I�     Y          �          
�  X�Y�     Z          �          
�  h�i�     [          �          
�  x�y�     \          �          
�  ����     ]          �          
�  ����     ^   |��.@�W�/�1��  
�  ����     _   |��.@�W�/�1��    @l��    Q     ��  h   h�
�  ���      �         @          
�  ���      +         @          
�  ` u!     ~          �          
�  x,yA     �          �          
�  �,�A               �          
�  �,�A     W          �          
�  �,�A     X         @            t�,    `     ��  ,   h�
�  P�Q      �         @          
�  0�1      P                     
�   %!     Q          �          
�  (,)A     R         @          
�  8,9A     S          �          
�  H,IA     T          �          
�  X,YA     U         @            $\,    h     ��  ,   ��  CClock
�  8�9�     P                       4�<�    q   ����     ��  CLED_G
�  8� M�      9          �          
�  d� y�      M                       L� d�     t   ��      r�
�  8� M�      :          �          
�  d� y�      M                       L� d�     w   ��      r�
�  8x My      ;          �          
�  dx yy      M                       Ll d�     z   ��      r�
�  8X MY      <          �          
�  dX yY      M                       LL dl     }   ��      r�
�  88 M9      =   B��� @ �:�?  
�  d8 y9      M            �:��    L, dL     � 
 ��      r�
�  8 M      >          �          
�  d y      M                       L d,     �   ��      ��  � �     220        �k@      �?   
�  � �      6 	        �          
�  �( �)      5 	 �v��D/@'�:�?  
�  �8 �9      4 	        �          
�  �H �I      3 	        �          
�  �X �Y      2 	        �          
�  �h �i      1 	        �          
�  �x �y      0 	        �          
�  �� ��      / 	        �          
�  �� ��      7          �          
�  �x �y      8          �          
�  �h �i      9          �          
�  �X �Y      :          �          
�  �H �I      ;          �          
�  �8 �9      <          �          
�  �( �)      =   B��� @'�:��  
�  � �      >          �            � ��      �     �� v   ��  CCounter10B
�  H8 ]9      �         @          
�  HH ]I      +         @          
�  HX ]Y      8          �          
�  h� i�      -          �          
�  x� y�      .          �          
�  �� ��      /          �          
�  �x �y      0          �          
�  �h �i      1          �          
�  �X �Y      2          �          
�  �H �I      3          �          
�  �8 �9      4          �          
�  �( �)      5   �v��D/@@�:��  
�  � �      6          �            \ ��      �     ��( T     H � H �     ���  CWire  HX I�       8 ��  H� 	�      8 ��  x 	�       8 ��  �x 	y      8 ��  � �� 	      � ���� 
 CCrossOver  � �� �        � �	�     � ����  � �� �        � �� 	      � ��  �	)      � ��  � `� i      � ����  � T� \        � P� a      � ����  � \� d        � `� a     � ����  � T� \        � H� a      � ����  � \� d      ��  � T� \        � P� i      � ����  � T� \      ��  � T� \      ��  � T� \      ��  � T� \      ��  � T� \      ��  � T� \        � XAY     � ��  � H� I     � ��  � 0� I      � ����  � T� \        � P� i      � ��  � ��     � ��  �  	     � ��  � 	     � ��  � �� !      � ��  � ��       | ��  � ��       � ��  � �� 	      } ��  �  � !     � ��  � � A      | ��  � � Q      � ��  x y a      } ��  � �� �     � ��  � ���     � ����  � T� \        � P� i      � ��  � P� Q     � ��  � �� Q      � ��  � h� i     � ����  ^ddl      ��  ^\dd        `Xaq      � ����  nTt\      ��  ~T�\      ��  �T�\      ��  �T�\        `X�Y     � ����  ^ddl      ��  ~d�l      ��  ndtl        Hh�i     � ����  ^\dd      ��  n\td        P`�a     � ����  ����        ���Y      � ��  ����     � ����  �T�\        �P�q      � ����  ����      ��  ����        x���     � ��  ����     � ��  P8Qa      � ��  HHIi      � ��  Ppaq     � ����  ����        ���	      � ��  x�y	      � ��  ���	      � ��  � �      | ��  � �      � ����  � T� \        � P� i      � ��  � X� i      � ��  @XAq      � ��  � PQ     � ��  � ��       � ��  �Q      � ��  � @	A     � ��  � �� 	      � ��   	A      � ��   1      � ��  � 01     � ��  �  � 1      � ��  � 0� 1     � ��  � @� A     | ��  � P� Q     � ��  x `� a     } ��  x � 	     } ��  ()i      G ��  @�A      G ��  (A     G ��  (hIi     G ��  P�Q      F ��  0Q     F ��  8 a!     E ��  01Y      F ��  0XIY     F ��  `�a!      E ��  8 9I      E ��  8HII     E ��  @8I9     D ��  @(A9      D ��  @(q)     D ��  p�q)      D ��  �8�9     C ��  ��9      C ��  ��I      B ��  ��     C ��  ���      C ��  �H�I     B ����  ���        ���Y      A ��  ��	     B ��  ���	      B ����  ����        ����     A ��  �X�Y     A ��  �h�q      � ��  H8Q9     � ����  ~d�l        �`�q      � ��  X(Y1      � ��  (Y)     � ����  nTt\      ��  n\td      ��  ndtl        pPqq      � ����  ~T�\        �P�a      � ����  �T�\        �P�i      � ��  (	A      � ����  ����        �P�      � ��   �!	      � ����  >�D�         �a�     � ��  `�a)      � ����  >�D�        @�A	      � ��  @���     � ��  ��A�     � ����  ��        ���I      � ��  �H	I     � ����  ��        �	     � ����  T\      ��  \d        H	i      � ��  �h	i     � ����  T\      ��  FTL\      ��  6T<\      ��  &T,\      ��  T\        �X�Y     � ��  `(aA      � ��  �Y�     � ��   �	�     � ����  ��        �	Y      � ����  ��      ��  ����        ��A�     ~ ����  �T�\      ��  �T�\      ��  �T�\      ��  �T�\        �X	Y     � ��  ���     � ����  �T�\        �P�q      � ����  �T�\        �P�i      � ����  �T�\        �P�a      � ����  �T�\      ��  �\�d      ��  �d�l        �P�q      � ����  �\�d      ��  �d�l        �X�q      � ��  �p�q     � ����  �\�d      ��  �\�d        �`�a     � ��  �8�a      � ����  �d�l      ��  �d�l      ��  �d�l        �h�i     � ��  `(�)     � ��  �(�1      � ����  �d�l        �`�q      � ��  �8�9     � ��  �H�i      � ��  �h�q      � ��  ���	      ~ ����  ����        ���	      � ��   `�      � ��   8 a      � ��  �XY     � ��  ���     � ��  ���	      � ��  �	     � ��  �Y      � ��  �HI     � ��  ���      � ��  �	     � ��  I      � ��  	9      � ��  �8	9     � ��  ���)      � ��  �(�)     � ��  �(�9      � ��  �8�9     � ��  �H�I     � ��  � �I      � ��  ���!      � ��  �X�Y     � ��  ��Y      � ��  � �!     � ��  ��     � ��  ���      � ��  �h�i     � ��  ��     � ��  ���      � ��  ��i      � ��  ��	     � ��  ��a      � ��  �`�a     � ��  ��Q      � ��  �P�Q     � ��  ��A      � ��  �@�A     � ��  �0�1     � ��  � �1      � ��  � !     � ��  H0Y1     � ��  XY1      � ��  ` aA      � ��  (�)	      � ��  H@aA     � ��  h�iQ      � ��  8�9      � ��  HPiQ     � ��  �X�q      � ��  (`)i      � ����  \d      ��  T\        Pi      � ����  �\�d        �X�i      � ����  &T,\        (P)a      � ����  \d      ��  �\�d      ��  \d        �`)a     � ��  �P�a      � ��  �P�Q     � ��  �H�Q      � ��   1      � ��  8`9i      � ����  F\Ld      ��  FTL\        HPIi      � ����  N�T�        H�i�     � ����  N�T        8 a     � ����  NT        (Y	     � ����  6T<\        8P9a      � ����  F\Ld        8`Qa     � ����  NT      ��  N�T      ��  N�T�        P`Q      � ��  ��     � ��  �	     � ��   Q     � ��    !      � ����  �        �!      � ����  �        �	      � ����  ���        ���      � ����  ���        ���	      � ����  ���      ��  ���      ��  ���      ��  �      ��  �        � !     � ��  �P�Q     � ��  �H�Q      � ��  889A      W ��  @9A     W ��  @�      W ����  F�L�      ��  V�\�      ��  f�l�      ��  v�|�        ���     W ����  F�L�        H�I�      v ����  V�\�        X�Y      u ����  f�l�        h�i	      t ����  v�|�        x�y      s ��  ���      W ��  � �     W ��  @i	     t ��  8 Y     u ����  ����      ��  ����      ��  ����        �P�      W ����  �L�T        �P�Q     W ����  �D�L        �@�Q      W ����  ����        ����     z ����  ����        ����     y ����  ����        ����     x ����  �L�T      ��  �D�L        �@�Y      X ��  �P�Y      W ��  `�a!      ~ ����  V�\�        @�a�     ~ ����  V�\�        X�YA      � ��  H8IA       ��  @@IA      ��  @@AQ       ����  FLLT      ��  fLlT      ��  vL|T        @P�Q      ����  �D�L        �@�Q       ����  FLLT        HHIY      M ����  fLlT      ��  fDlL        h@iY      � ����  vL|T      ��  vD|L        x@yY      � ��  �P�Y       ����  fDlL      ��  �D�L      ��  �D�L      ��  �D�L      ��  vD|L        HH�I     M ����  ~���        ����      + ��  ����      � ��  XXiY     � ��  � �     R ��  � �A      R ����  �<�D        �@)A     R ��  �`a     � ����  ����        ���     U ����  �<�D      ��  ����      ��  ����        ���I      M ��  ����     + ����  ����        ���A      + ��  �@�A     + ����  VL\T        XHYa      U ��  X@YI      U ����  fDlL        XHqI     U ����  fDlL        h�iQ      � ����  ��        ��      U ��  ���      U ��  �H�a      M ��  �@�A     x ��  ����      y ��  ���A      x ��  �0�1     y ��  ����      z ��  ���1      y ��  ���!      z ��  � �!     z ��  Hy     s ��  HI!      s ��  H Q!     s ��  @0Q1     t ��  @A1      t ��  8@QA     u ��  8 9A      u ��  0PQQ     v ��  0�1Q      v ��  0�I�     v ��  � �Y      i ��  `a     � ��  Pa      � ��  P�i�     � ��  P�Q�      � ����  VL\T      ��  FLLT      ��  6L<T      ��  &L,T        PiQ     � ����  FLLT        H@Ia      T ����  6L<T        8@9a      S ����  &L,T        (@)a      R ��  ���      i ��  � �     i ��  �XY     i ��  �		      j ��  �		     j ��  �     k ��  ��I      j ��  �HI     j ��  �      k ��  ��9      k ��  �89     k ��  �()     l ��  ��)      l ��  �)     l ��  (�)      l ��  X(i)     m ��  h i)      m ��  p�q9      n ��  8 i     m ��  8�9      m ��  X8q9     n ��  x�yI      o ��  H�q�     n ��  H�I�      n ��  X�y�     o ��  XHyI     o ����  ~���        X���     � ����  6�<�        �q�     U ����  6�<�      ��  ����      ��  ��      ��  ����        ��Q�     � ����  6�<�      ��  6�<�        8�9�      P ��  0�9�     P ��  p�qI      U ��  �� ��      M ��  �� ��       M ��  x� ��      M ��  �x ��       M ��  x� ��      M ��  �X �y       M ��  xx �y      M ��  �8 �Y       M ��  xX �Y      M ��  � �9       M ��  x8 �9      M ��  x �      M ��  � 9�      9 ��  h �       9 ��  �h i      9 ��   X !�       : ��   � 9�      : ��  �X !Y      : ��  (H )y       ; ��  (x 9y      ; ��  �H )I      ; ��  08 1Y       < ��  0X 9Y      < ��  �8 19      < ��  8( 99       = ��  �( 9)      = ��  � 9      > ��  X@iA     � ��   8 I9      � ��   ���     M ��   �!�      M ��  ��!�     M ��  p���     + ��  pq�      + ��  q     + ��  H       + ��  H II      +   H � H �     �  H � H �       H � H �      2   g   f   e   d   c   b   a            �  �  �  �       �" " # 	# $ 
$ % % & & , ' '   ( ( �) ) * * , & , . . / / 0 0 1 1 2 2  3 3   4 4 )5 5 "6 6 9 X 9 : W : ; V ; < U < = T = > S > ? R ? @   @ A A   B B C C D D E E F F !G G &H H 'K �K L *L M ,M N 0N O �O P �P Q �Q R R ? S S > T T = U U < V V ; W W : X X 9 Z �Z [ �[ \ �\ ] �] ^ �^ _ �_ ` �` a a  b b  c c  d d  e e  f f  g g  j �j k �k l �l m m �n n �o o �p p �r �r s �s t .t u u 0v v 4w w 6x x �{ { �| | +} 8}   {� � z� R� � ~� � }� � w� � � f� � d� � b� � `� ?� � ;� � �� � � �� � �� � �� � �� �� � �� � �� � �� � K� � K� � �� � � � � � � � � � � � � � � � � � � � � � � `� � |� � x� � f� � m� � m� � �� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �   � � �   � � �� � �� � �� � �� � �� � �� � �� �� � �� � �� � �� � � � � �   � � �� � �� � �� � � � �� � �� � �� � �� � � � � �   � � �� � �� � �� � � � � � � � � � � � � � � � � � � � � �   � � �   � � �� � �� � �� � �� � �� � �� � �� � � � � �� � �� F� � � �� � � � � � � �   � � � � � � 1 * -E;^]	\	
[
ZYX    ����KHQRTV"  GJ  N""$$4&t&'s'(p()k)** ++  ,,�--}..x1O12N23M34L45K56J67I78  899  ::i;;l<<q==w>>|??�@@�B<BCcCDeDEgEF[FGZGHFHII7JJ6KK5LL4MM3NN2OO1QQRRS"STTU,UV,VWWXXYYZZ[[
\\	]]^^`+`a)abbccddee ffh]hi�ij  jkkgllemmcnn>qq�t�tuu�w�wxx�z�z{{�}�}~~���������������������������������������  ��������������������������������  ��  ���������������������������������k �������j �/�\ ��n �������������m ] ����������������l ���p Z    � � � ��	�
�������^ ����_ ������O �1�5�7�������-�3�*���2�,��������x K �������B+�{ �P ����r �s �� ������o [ �` �Q (  ���)  ���* �" �# �$ �% ��B 1 C 0 D / . E 6  %"!F  5 #�')&G %':H #4 #6L | �,�4M /t 8.0�0�0�u N 4�v �6�w ��} 9(��<� <@;><R?=B� ?~CACG�ECHFD��HMH�E� � HLIL�L�L�L���v� T�UUXSZWVW}� ZgZeZcZajUAT`^� � b]� rd\� nf[fpfu� � jojsZ� � jnknhqxznrlryri{|>wv� xtd� � q rb� W� ~Y_� �_�1� �� �� ������ �� �������� �� ������� �� ��� ��� ������� ��� ��� ��������� ���� ���� �� ����� ������ �� ���� �� �L� �� ���Q� � ��L� �P� ��J����������� �F� �� ���N� � ��� ����������O� ������������������������ ���� ���� ���� ��$��������9�9�� �� �����������������X��������O����S�U�������	� &e��KM�HL�I�%fQ RbW���  "'d#W$�U(cTS##
###!F)��a�`V.-//5.k� �26EC40434��#)99�8;9<_>Bn??B<�A@\^C��224HIGLJN MP�OQPS�RU�TWXVW�jkGF^Z�A\h^=^d^f^h[Ac`mCealDgb/E:jYiY);molrqmpo(<nnsr'u&vtuw=v.y{x}|y>{-z���z?@~,~�*S+��C����:�D�7�]����q�i��?����u���x���{���~��������t�������w�����z�����}��������������$��8�������� �          �$s�        @     +        @            @    "V  (      �                
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 