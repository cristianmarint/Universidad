��  CCircuit��  CSerializeHack           ��  CPart              ���  CAND�� 	 CTerminal  ��	               �          
�  ��               �          
�  ��               �            ��           ��    �� 	 CInverter
�  P(e)              @          
�  |(�)               �            d|4           ��    ��  CNOR
�  @� U�               @          
�  @U	              @          
�  l �               �            T� l           ��    ��  CLED_G
�  ����       	        �          
�  ����                            ���         ��      �� 	 CResistor��  CValue  �q�    330          �t@      �?   
�  �X�m                �          
�  ����               �            �l��         ��      ��  CLED_Y
�   h!}       	 �y����?�kl�ʣ�?  
�   �!�                �kl�ʣ��    |4�     #  	 ��      �
�  phq}       	 ����� @�}"T�?  
�  p�q�                �}"T��    d|��     &   ��      ��  �AO    330          �t@      �?   
�   (!=               @�kl�ʣ�?  
�   T!i        �y����?�kl�ʣ��    <$T     *    ��      ��  KAkO    330          �t@      �?   
�  p(q=               @�}"T�?  
�  pTqi        ����� @�}"T��    l<tT     .    ��      ��  CBattery�  � � � �     5V(          @      �? V 
�  � � � �                @�tG}U��  
�  � � � �                 �tG}U�?    � � � �      3    ��      ��  CSPST��  CToggle  x� ��      6   
�  p� q�               @�}"T��  
�  p� q�                @�}"T�?    l� t�     9     ��    5�7�  (� H�      ;   
�   � !�               @�kl�ʣ��  
�   � !�                @�kl�ʣ�?    � $�     =     ��    ��  CEarth
�  � p� �                       ��    � �� �     A    ��                    ���  CWire  �X�Y      C�  ��Y       C�  PQ)       C��� 
 CCrossOver  $        pQ      C�  pq       C�H�  $      H�  $         � !)       C�  pq)       C�  ��)       C�  ��	      C�  � �	       C�  p� q	       C�H�  $        pA	      C�  @� A�        C�   � A�       C�   � !�        C�   �!�       C�   �!�       C�   ���      C�  p�!�      C�  � � q�       C�  � � � a       C�  �q�      C�  p�q�       C�  � `� q       C�  � `	a      C�  `	�       C�  p� !�                     �                             P   O    E  F    O  U   S    Q       Z  D       # + # $ $ Y & / & ' ' _ * K * + + # . N . / / & 3 \ 3 4 4 ] 9 9 R : c : = = W > c > A ` A E   D G  G L N F R G K I K T W * J .   Q   P 9 S S M J  V  K U = V Y [ $ Z X  ^ X 3 : 4 a b _ ' [ ] A ` b a ^ \ >             �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 