��  CCircuit��  CSerializeHack           ��  CPart    0   0     ���  CECapacitor��  CValue  ���    100�F(    -C��6?      �?�F �� 	 CTerminal  ��         �H���?ʒ)d,`�  �  �                ʒ)d,`?    ��        ��      q��gC��>��  CLED�  ����       	 �g:.��? X�F�Ċ?  �  ����                 X�F�Ċ�    ����       
 ��      ��  p�q�       	 �g:.��? X�F�Ċ?  �  p�q�                 X�F�Ċ�    d���       
 ��      ��  P�Q�       	        �          �  P�Q�                            D�d�         ��      ��  0�1�       	        �          �  0�1�                            $�D�         ��      �� 
 CResistors
�  	i)w    220          �k@      �?   �  �P�e                �          �  �P�e      
   �o�� @#X�F�Ċ?  �  �P�e                �          �  pPqe         �o�� @#X�F�Ċ?  �  `Pae                �          �  PPQe                �          �  @PAe                �          �  0P1e                �          �  0|1�               �          �  @|A�               �          �  P|Q�               �          �  `|a�               �          �  p|q�        �g:.��?#X�F�Ċ�  �  �|��               �          �  �|��        �g:.��?#X�F�Ċ�  �  �|��               �            *d�|          �� v   �� 	 CPushMake��  CKey  �Z�v      0   �  �t��              @          �  �H�]       	        �            �\�t    3      ��    �� 
 CCounter16�  ��	              @          �  �(�)               �          �  �4�I               �          �  �0�1               �          �  � �!               �          �  ��        �o�� @ X�F�Ċ�  �  � �     
   �o�� @ X�F�Ċ�    �� �4     7      ��  ,   ��  CBattery
�  !3/    5V(          @      �? V �  @A               @z(=e��  �  @4AI                z(=e�?    4L4     A    ��      ��  CEarth�  @HA]       	         z(=e��    3\Kd     E    ��      ��  CSPST��  CToggle  ��0     G   �  ��	              @z(=e�?  �  ��	              @z(=e��    ��     J     ��    �� 	 CResistor
�  ���    220          �k@      �?   �  ��       	        �          �  �                            ��     O    ��      ��  CLED_G�  ��                �          �  ��               �            �$�     S    ��      C��  (=                 �J��g�?    <D     V    ��      ��  C555�  �(�=               @N贁Nk?  �  �(�=               @          �  �@�A     	   �H���?��8��J�?  �  �P�Q        �H���?          �  �`�a        �H���?          �  �d�y                ao9 ?��  �  �d�y        ������
@       �  �  �P�Q               �            �<�d     Y    ��   (   �� 
 CVResistor��  CSlider   t/�     
�  ���    0k     F]t�1�@        k 
   e �  h}      	 	 �H���?Ȓ)d,`�  �  ��        �H���?Ȓ)d,`?    |�     f    ��      L�
�  �AO    470          `}@      �?   �  (=               @<s���?�?  �  Ti     	   �H���?<s���?��    <T     j    ��          0   0     ���  CWire  Pq      m�  p�      m�  ���       m�  0Q      m�  p�q       m�  1      m�  P�Q       m�  �      m�  0�1       m�          m�  �i	      m�  �	      m��� 
 CCrossOver  fLlT        P�Q      m�  � �Q      
 m�  � �     
 m�  pqQ       m�  �q      m�  � Q!      m�  P QQ       m�  001Q       m�  �011      m�  �(�Q       m�{�  fLlT        hi�       m�  h���      m�  h�	      m�  �      m�  �x�       m�  �	      m�  @�	      m�  )       m�         m�  P�       m�  �PQ      m�  p`q�       m�  pPqa       m�  p`�a      m�  hai     	 m�  ��       m�  ��       m�  �q�      m�  pP�Q      m�  `@ai      	 m�  `@�A     	 m�  ��)       m�  ��	      m�  ��)       m�  )           0   0     �    0   0         0   0      �    �  -    p  +    r  )    t  '    v       }   !   ! "  " #   # $ � $ %   % & � & ' '  ( (   ) )  * *   + +  , ,   - -  . .   3 3 � 4 9 4 7 � 7 8 � 8 9 9 4 : : � ; ; � < < � = = ~ A � A B B E E B E J � J K K � O T O P P w S � S T T O V � V Y � Y Z � Z [ � [ \ � \ ] � ] ^ ^ � _ _   ` ` � f k f g g � j � j k k � q r n p  o s t  o u v  n � w  q P s � � � � z � � � ~   = } � " <  ; � � $ � & : � 8 z � | � � � 3 x 7 � � ^ u K y A J � V  � � S ` z � � � � � ] f � �  g � � � � \ � � � [ � Y � x y Z � j            �$s�        @     +        @            @    "V  (      �P                
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 