��  CCircuit��  CSerializeHack           ��  CPart              ��� 	 CInverter�� 	 CTerminal  � �               �          
�  �               @            �� �           ��    ��  COR
�  � %�               @          
�   %      	       @          
�  <� Q�         ���P�p@����\*��    $� <           ��    �
�  �� ��                �          
�  � !�               @            �� �            ��    �
�  �� ��                �          
�  �� ��               @          
�  �� 	�               @            �� ��            ��    ��  CLED_G
�  � �         �٭$M� @����\*�?  
�  �,�A                ����\*��    ��,        ��      �� 	 CResistor��  CValue  ����    330          �t@      �?   
�  �x��         ���P�p@����\*�?  
�  ����        �٭$M� @����\*��    ����     !    ��      ��  CSPST��  CToggle  �x ��       $   
�  �� ��                �          
�  �h �}                @            �| ��     '      ��    #�%�  �x �       )   
�  �� ��                �          
�  �h �}                @            �| ��     +      ��    #�%�  p 0�       -   
�  � 	�                �          
�  ` 	u                @            t �     /      ��    ��  CBattery�   � 3 �     5V(          @      �? V 
�  @ � A �                @          
�  @ A                             4 � L      4    ��      ��  CLED_Y
�  ��      	          �          
�  �4�I                            ��4     8    ��      6�
�  � �                �          
�  �,�A                            ��,     ;    ��      6�
�   	                �          
�  ,	A                            � ,     >    ��      ��  ����    330          �t@      �?   
�  �x��                �          
�  ����     	          �            ����     B    ��      ��  ����    330          �t@      �?   
�  �x��                �          
�  ����               �            ����     F    ��      ��  � ��    330          �t@      �?   
�  x	�                �          
�  �	�               �            ��     J    ��      ��  CEarth
�  @ �A �                 ����\*�?    3 �K �     N    ��                    ���  CWire  � 	y       P�  � 	�        P��� 
 CCrossOver  �� ��       T�  �� ��         � ��       P�  �� ��        P�  �� �y       P�  P� ��       P�  � �	       P�  ��	      P�T�  �� ��       T�  �� ��         �� �	       P�  ��y       P�  � �        P�  � �       P�T�  �� ��          � ��       P�T�  �� ��         �� ��        P�  �� �y       P�   	a        P�  � �i        P�  ����      P�  ����      P�  �@��       P�  ���       P�  � �i        P�  � �       P�   �       P�  @  	       P�  @  A �        P�  X �q �      P�  @ �Y �      P�  X �Y �       P�  @ �Y �      P�  @ A �       P�  @ �A �       P�  ���      P�  �H��       P�  @	�       P�  �@��       P�  p �q �       P�  p �	�      P�  ���	      	 P�  ���       P�  �	                     �                             Z      `       Y  f    b  S   W    a  l    k ! X ! " " l ' ' \ ( m ( + + d , h , / / R 0 g 0 4 q 4 5 5 v 8 ~ 8 9 9 y ;  ; < < { > � > ? ? z B _ B C C ~ F f F G G  J Q J K K � N w N R J / S S e S ] Q   b Y !  X  [ _ Z \ V \ c ' [ \ B a   ` b ^  W d U +  d F p 0 o , x y i k  j "  n ( h m g n q o p 4 s | w t u r v t 5 u s N z { 9 j ? } < i r } | x C 8 G ; K >             �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 