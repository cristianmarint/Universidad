��  CCircuit��  CSerializeHack           ��  CPart              ���  CAND�� 	 CTerminal  �(�)              @          
�  �8�9              @          
�  �0�1        ���P�p@����\*��    �$�<           ��    �
�  @� U�               @          
�  @ U              @          
�  l� ��               @            T� l           ��    ��  CLED_G
�  � �         �٭$M� @����\*�?  
�  �,�A                ����\*��    ��,        ��      �� 	 CResistor��  CValue  ����    330          �t@      �?   
�  �x��         ���P�p@����\*�?  
�  ����        �٭$M� @����\*��    ����         ��      �� 	 CInverter
�   859               �          
�  L8a9              @            4,LD           ��    �
�  ��	               �          
�  !	              @            ��      !      ��    �
�  �� ��                �          
�  �� ��               @            �� ��      $      ��    ��  COR
�  �� �                �          
�  �� �       	       @          
�  $� 9�               @            � $�      (      ��    ��  CSPST��  CToggle  �x ��       ,   
�  �� ��                �          
�  �h �}                @            �| ��     /      ��    +�-�  �x �       1   
�  �� ��                �          
�  �h �}                @            �| ��     3      ��    +�-�  p 0�       5   
�  � 	�                �          
�  ` 	u                @            t �     7      ��    ��  CBattery�   � 3 �     5V(          @      �? V 
�  @ � A �                @          
�  @ A                             4 � L      <    ��      ��  CLED_Y
�  ��      	          �          
�  �4�I                            ��4     @    ��      >�
�  � �                �          
�  �,�A                            ��,     C    ��      >�
�   	                �          
�  ,	A                            � ,     F    ��      ��  ����    330          �t@      �?   
�  �x��                �          
�  ����     	          �            ����     J    ��      ��  ����    330          �t@      �?   
�  �x��                �          
�  ����               �            ����     N    ��      ��  � ��    330          �t@      �?   
�  x	�                �          
�  �	�               �            ��     R    ��      ��  CEarth
�  @ �A �                 ����\*�?    3 �K �     V    ��                    ���  CWire  �x�y      X�  �0�y       X�  �� �)       X�  `8�9      X�  8� 9�        X�  @ A	       X�   A	      X�  8� A�       X�  ����      X�  ����      X�  �@��       X�  ���       X�  �8�y       X��� 
 CCrossOver  �� ��       g�  �� ��       g�  ��        �� �9       X�  �8!9      X�   	a        X�  � �i        X�  ��y       X�g�  �� ��       g�  �� ��         �� �	       X�g�  ��        ��	      X�  � 	y       X�  � 	�        X�g�  �� ��       g�  �� ��         � ��       X�  � 	�        X�g�  �� ��       g�  �� ��         � ��       X�  � �i        X�  � �       X�   �       X�  @  	       X�  @  A �        X�  X �q �      X�  @ �Y �      X�  X �Y �       X�  @ �Y �      X�  @ A �       X�  @ �A �       X�  ���      X�  �H��       X�  @	�       X�  �@��       X�  p �q �       X�  p �	�      X�  ���	      	 X�  ���       X�  �	                     �                             [   \    Z  `   ^    [  d    c  Y    d  k    \ ! r ! " " _ $ v $ % % ) ( z ( ) % ) * * ] / / f 0 } 0 3 3 o 4 m 4 7 7 y 8 l 8 < � < = = � @ � @ A A � C � C D D � F � F G G � J e J K K � N n N O O � R t R S S � V � V  Z  Y     * `  _ " ^ ]  � � a c  b   f J f | f x f s / k e  � 8  4 o N o { o w 3 r r j n ! u R y v v q v i t $ 7 z z p z h u ( ~ 0 m } l ~ �  � < � � � � � � � � = � � V � � A b G � D a � � � � K @ O C S F             �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 