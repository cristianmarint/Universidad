��  CCircuit��  CSerializeHack           ��  CPart    0   0     ���  CLED_G�� 	 CTerminal  � �!     1          �          
�  � �!                            ��4        ��      �
�  �@�A     2          �          
�  �@�A                            �4�T        ��      �
�  �`�a     3          �          
�  �`�a                            �T�t        ��      �
�  ����     4          �          
�  ����                            �t��        ��      �
�  ����     5          �          
�  ����                            ����        ��      �
�  � �     0          �          
�  � �                            �� �        ��      �
�  �� ��      /          �          
�  �� ��                             �� ��         ��      �
�  �� ��      .   B��� @ �:�?  
�  �� ��                  �:��    �� ��        
 ��      �
�  �� ��      -          �          
�  �� ��                             �� ��     #    ��      �
�  �� ��      ,          �          
�  �� ��                             �t ��     &    ��      �� 
 CResistors��  CValue  �    220        �k@      �?   
�  � �!     '          �          
�  �0�1     (          �          
�  �@�A     6          �          
�  �P�Q     7          �          
�  �`�a     8          �          
�  �p�q     9          �          
�  ����     :          �          
�  ����     ;          �          
�  �)�     <          �          
�  �)�     =          �          
�  p)q     +          �          
�  `)a     	          �          
�  P)Q               �          
�  @)A     *          �          
�  0)1     5          �          
�   )!     4          �            ��     ,      �� v   (�*�  �n |     220        �k@      �?   
�  �� ��       	        �          
�  �� ��        	        �          
�  �� ��      ! 	 �v��D/@'�:�?  
�  �� ��      " 	        �          
�  �� ��      # 	        �          
�  �� ��      $ 	        �          
�  �� ��      % 	        �          
�  �� ��      & 	        �          
�  � )�      3          �          
�  � )�      2          �          
�  � )�      1          �          
�  � )�      0          �          
�  � )�      /          �          
�  � )�      .   B��� @'�:��  
�  � )�      -          �          
�  � )�      ,          �            �| �      >      �� v   ��  CCounter10B
�  �� ��               @          
�  �� ��                �          
�  �� ��      )          �          
�  �� �	     (          �          
�  �� �	     '          �          
�  �� ��      &          �          
�  �� ��      %          �          
�  �� ��      $          �          
�  �� ��      #          �          
�  �� ��      "          �          
�  �� ��      !   �v��D/@@�:��  
�  �� ��                 �          
�  �� ��                �            �| ��      P      ��( T   ��  CAND
�  ����               �          
�  ����               �          
�  ����                �            |���    _      ��    ��  CSevenSegmentDisplay
�  xP�Q        �i�n� @ W�/�1�?  
�  x`�a               �          
�  xp�q        �i�n� @ W�/�1�?  
�  x���        �i�n� @ W�/�1�?  
�  ����                �l��~��  
�  ����               �          
�  �p�q               �          
�  �`�a        �i�n� @ W�/�1�?  
�  �P�Q        �i�n� @ W�/�1�?    �L��     d 	     ��0 <             (�*�  ��    220        �k@      �?   
�  ��      	        �          
�  � �!      	 |��.@�W�/�1�?  
�  �0�1      	 |��.@�W�/�1�?  
�  �@�A      	 |��.@�W�/�1�?  
�  �P�Q      	        �          
�  �`�a      	 |��.@�W�/�1�?  
�  �p�q      	 |��.@�W�/�1�?  
�  ����               �          
�  �)�               �          
�  p)q        �i�n� @�W�/�1��  
�  `)a        �i�n� @�W�/�1��  
�  P)Q               �          
�  @)A        �i�n� @�W�/�1��  
�  0)1        �i�n� @�W�/�1��  
�   )!        �i�n� @�W�/�1��  
�  )               �            ��     o      �� v   ��  C4511
�  ��               �          
�  � �!     
         @          
�  �0�1               �          
�  �@�A               �          
�  �P�Q              @          
�  �`�a              @          
�  �p�q              @          
�  �p�q        |��.@�W�/�1��  
�  �`�a        |��.@�W�/�1��  
�  �P�Q               �          
�  �@�A        |��.@�W�/�1��  
�  �0�1        |��.@�W�/�1��  
�  � �!        |��.@�W�/�1��  
�  ��               �            ��x     �      ��  h   �� 	 CPushMake��  CKey  Rjv�      �   
�  H�I�              @          
�  HXIm       	        �            @lL�    �      ��    �� 
 CCounter10
�   5              @          
�   859              @          
�  HDIY               �          
�  T@iA               �          
�  T0i1               �          
�  T i!     
         @          
�  Ti               �            4TD     �      ��  ,   ��  CSPST��  CToggle  �  � @     �   
�  x �       	       @          
�  � �               @            � �      �     ��    �� 	 CVoltRail*�  3 [     5V(          @      �? V 
�  d y               @            \ d      �    ����     ��  CClock
�  L pa q              @            4 lL t     �    ����     ��  CEarth
�  ����       	         @y����?    ����     �    ��          0   0     ���  CWire   � ��       ��   � !       ��  !      ��  �@�A      ��  h@�A      ���� 
 CCrossOver  �,�4      ��  ��$      ��  ��        ���A       ����  �,�4        h0�1      ����  ��$        h �!     
 ����  ��        ��      ��  h�      ��  ���       ��  �� ��       ��  �� ��       ��  �0�1     ( ��  ��1      ( ��  � �!     ' ��  ��!      ' ��  �	�       ��  �	�       ��  ��	�      ��  `	�       ��  ��	�      ��  @	a       ��  �`	a      ��   	A       ��  �@	A      ��   	!       ��  � 	!      ��  � 	       ��  � 	      ��  � 	�        ��  �� 	�       ��  � 	�        ��  �� 	�       ��  � 	�        ��  �� 	�       ��  ��	�      ��  �� 	�       ��  H���     5 ��  H0I�      5 ��  (0I1     5 ��  P Q�      4 ��  X� Ya      3 ��  P���     4 ��  ( Q!     4 ��  X`�a     3 ��  (� Y�      3 ��  `� aA      2 ��  `@�A     2 ��  (� a�      2 ��  h �!     1 ��  h� i!      1 ��  (� i�      1 ��  p� q      0 ��  p �     0 ��  (� q�      0 ��  x� y�       / ��  x� ��      / ��  (� y�      / ��  �� ��       . ��  �� ��      . ��  (� ��      . ��  �� ��       - ��  (� ��      - ��  (� ��      , ����  � \� d      ��  \d        � `!a      ��  �p��       ��  �p�q      ��  �`�a      ��  �P�a       ��  �P�Q      ��  �`��       ��  `pa�       ��  `�y�      ��  hpyq      ��  h`iq       ��  p`ya      ��  pPqa       ��  (PqQ      ��  x@yQ       ��  (@yA      ��  �p�q      ��  ��q       ��  (�      ��  � �a       ��  ( �!      ��  �`�a      ��  �0�Q       ��  (0�1      ��  � 	      ��  � `� �       ��  ` p� q      ��  � 8� q       ����  � 4� <      ��  � \� d        � � �       ����  4<      ��  \d        	�       ��   8!a       ����  4<      ��  � 4� <        � 8!9      ��  � �       ��  (`ia      ��  (paq      ��  � ���      ��  � ���      ��  �I�          0   0     �    0   0         0   0      �    �  �    �  �    �  �    �  �    �  �    �  �    �   �   ! ! � # � # $ $ � & � & ' ' � , � , - � - .   . /   / 0   0 1   1 2   2 3   3 4 4   5 5   6 6   7 7   8 8   9 9   : : � ; ; � > \ > ? [ ? @ Z @ A Y A B X B C W C D V D E U E F F � G G � H H � I I � J J � K K � L L � M M � P � P Q � Q R   R S S � T T � U U E V V D W W C X X B Y Y A Z Z @ [ [ ? \ \ > _ _ � ` ` � a � a d d e e f f g g h h � i i   j j 
k k l l o � o p � p q � q r � r s � s t � t u � u v   v w w   x x "y y !z z { { 	| | } } ~ ~ � � � � � � � � � � � � � � � � � � � � � � � u � � t � � s � � r � � q � � p � � o � � %� � � � � � � � � � � � � � � � � � � � � � � � � � � �  � � � � � � � � � P � � � � � � � � � � � � � ` � � � � � � � � � � � � � � � _ � � Q � a � - S � � , T � � � � �  � � �  � � �  � � �  � � �  � � �  � � �  � � � ! � � � $ � h � ' � �  � � : � � � � � �  ; � �  F � � � �  G � �  � � H � � � �  I � � � �  J � � � �   K � � # L � M & � � � #� �  � � � � � � $"g f !e z 	d { j 
~ } k l | � #� �  $� � %� � � y x �  �  >          �$s�        @     +        @            @    "V  (      �P                
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 