��  CCircuit��  CSerializeHack           ��  CPart    0   0     ���  CECapacitor��  CValue  ���    100�F(    -C��6?      �?�F �� 	 CTerminal  ��         �7�@ �t5�?  �  �                 �t5��    ��        ��      �D���+?��  CBattery
�  !3/    5V(          @      �? V �  @A               @����7��  �  @4AI                ����7�?    4L4         ��      ��  CEarth�  @HA]       	         ����7��    3\Kd         ��      ��  CSPST��  CToggle  ��0        �  ��	              @����7�?  �  ��	              @����7��    ��          ��    �� 	 CResistor
�  ���    220          �k@      �?   �  ��       	 �P��@9 @Aj~�?  �  �                9 @Aj~��    ��          ��      ��  CLED_G�  ��         </��`@ !@Aj~�?  �  ��        �P��@ !@Aj~��    �$�     $  
 ��      ��  (=                 �����7�?    <D     '    ��      ��  C555�  �(�=               @=W)�?  �  �(�=               @          �  �@�A     	   ���G��@          �  �P�Q        �7�@          �  �`�a        �7�@          �  �d�y                N贁Nk�  �  �d�y        ������
@       �  �  �P�Q        </��`@\@Aj~��    �<�d     *    ��   (   �� 
 CVResistor��  CSlider   t/�     
�  ���    50k     F]t�1�@�������?k 
   6 �  h}      	 	 ���G��@��t5�?  �  ��        �7�@��t5��    |�     7    ��      �
�  �AO    470          `}@      �?   �  (=               @�t5�?  �  Ti     	   ���G��@�t5��    <T     ;    ��          0   0     ���  CWire  �      >�  �      >�  �x�       >�  �	      >�  �	      >�  @�	      >�  )       >�         >�          >�  P�       >�  �PQ      >�  p`q�       >�  pPqa       >�  p`�a      >�  hai     	 >�  ��       >�  ��       >�  �q�      >�  pP�Q      >�  `@ai      	 >�  `@�A     	 >�  ��)       >�  ��	      >�  ��)       >�  )           0   0     �    0   0         0   0      N    F  D         D    C   %   ! ! G $ H $ % %   ' E ' * T * + V + , S , - Q - . L . / / A 0 0   1 1 I 7 < 7 8 8 O ; W ; < < M @ G E A / ? W U  B   F '  @ ! ? I $ 1 H K P Q L J . 7 R O  8 P N J K - S M R , U * V T B + C ;  
          �$s�        @     +        @            @    "V  (      �P                
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 