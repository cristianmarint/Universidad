��  CCircuit��  CSerializeHack           ��  CPart              ��� 	 CResistor��  CValue  K�k�    330          �t@      �?   �� 	 CTerminal  ppq�         ���P�p@����\*�?  �  p�q�        �٭$M� @����\*��    l�t�         ��      ��  CLED_G�  pq         �٭$M� @����\*�?  �  p4qI                ����\*��    d�4        ��      �� 	 CInverter�  P@eA     
          �          �  |@�A              @            d4|L           ��    ��  COR�  ((=)              @          �  (8=9              @          �  T0i1        ���P�p@����\*��    <$T<           ��    ��   -!               �          �  D Y!              @            ,D,           ��    ��  CAND�  ��	              @          �  ��              @          �  )              @            �     !      ��    ��  �� ��               @          �  �� ��               @          �  �� ��               @            �� ��      %      ��    ��  ��	               �          �  ��	              @            �� �     )      ��    ��  h� }�               @          �  h� }�               @          �  �� ��               @            |� ��      ,      ��    ��  � %�                �          �  <� Q�               @            $� <�      0      ��    ��  �� ��                �          �  � )�               @            �� �      3      ��    ��  CSPST��  CToggle  Xx x�       6   �  P� Q�      
          �          �  Ph Q}                @            L| T�     9      ��    5�7�  �x ��       ;   �  �� ��                �          �  �h �}                @            �| ��     =      ��    5�7�  �x �       ?   �  �� ��                �          �  �h �}                @            �| ��     A      ��    5�7�  p 0�       C   �  � 	�                �          �  ` 	u                @            t �     E      ��    ��  CBattery
�   � 3 �     5V(          @      �? V �  @ � A �                @          �  @ A                             4 � L      J    ��      ��  CLED_Y�  PQ                �          �  P4QI                            Dd4     N    ��      L��  ��      	          �          �  �4�I                            ��4     Q    ��      L��  � �                �          �  �,�A                            ��,     T    ��      L��   	                �          �  ,	A                            � ,     W    ��      �
�  +�K�    330          �t@      �?   �  PxQ�      
          �          �  P�Q�               �            L�T�     [    ��      �
�  ����    330          �t@      �?   �  �x��                �          �  ����     	          �            ����     _    ��      �
�  ����    330          �t@      �?   �  �x��                �          �  ����               �            ����     c    ��      �
�  � ��    330          �t@      �?   �  x	�                �          �  �	�               �            ��     g    ��      ��  CEarth�  @ �A �                 ����\*�?    3 �K �     k    ��                    ���  CWire  PHQ�       m�  P�q�      m�  pHq�       m�  p�q	       m�  p0qq       m�  h0q1      m��� 
 CCrossOver  N� T�       u�  �� ��       u�  �� ��         P� i�       m�   �       m�  (8)A       m�  �@)A      m�u�  N� T�       u�  N� T�       u�  NT      u�  NT$        P� QA      
 m�  P@Qy      
 m�   	a        m�  ())       m�  � �i        m�  ��!       m�u�  NT$      u�  ��$      u�  ��$        X �!      m�u�  ��$      u�  �� ��         �� �y       m�   !      m�  � 	!       m�   	y       m�  �� �	       m�  �� �	       m�u�  NT        ��	      m�  �� ��        m�u�  �� ��       u�  �� ��         �� �	       m�u�  ��$        ��y       m�  h� i�        m�u�  N� T�       u�  �� ��         (� i�       m�  � �       m�  � 	�        m�  �� ��       m�  �� ��        m�  P Qi        m�  � Q       m�  � �i        m�  � �       m�  @  	       m�  @  A �        m�  X �q �      m�  @ �Y �      m�  X �Y �       m�  @ �Y �      m�  @ A �       m�  @ �A �       m�  ����      m�  ��Q�      m�  ���      m�  �H��       m�  @	�       m�  �@��       m�  p �q �       m�  p �	�      m�  P�Q	       m�  ���	      	 m�  ���       m�  �	                     �                             r    q  q    p  �    {  �   z    s  �    � ! � ! " � " # # � % � % & � & ' ' � ) � ) * * � , � , - � - . . � 0 � 0 1 1 t 3 � 3 4 4 � 9 9 | : � : = = � > � > A A � B � B E E � F � F J � J K K � N � N O O n Q � Q R R � T � T U U � W � W X X � [ � [ \ \ � _ � _ ` ` � c � c d d � g � g h h � k � k O � n p  o   s   r t ~ t � t � 1 � � �  {  z | � | v | � | � 9  | [ � F #  y B " � � � � � � �  � � � � x � c �  � � � g ' ! & � �  * � . % � � � w = ) � � � _ - t � } � � 4 , � 0 E � � 3 A � � : � � � > � � � y � J � � � � � � � � K � � k � � � o � � R � X � U � � � � � \ N ` Q d T h W             �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 