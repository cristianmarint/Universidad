��  CCircuit��  CSerializeHack           ��  CPart�� 
 CTextLabel  � ��    Decodi.          �   �     ���  CCounter10B�� 	 CTerminal  (P =Q      S         @          �  (` =a      +         @          �  (p =q      >          �          �  H� I�      g          �          �  X� Y�      f          �          �  d� y�      {          �          �  d� y�      z          �          �  d� y�      y          �          �  dp yq      x          �          �  d` ya      w          �          �  dP yQ      v   �v��D/@@�:��  �  d@ yA      u          �          �  d0 y1      t          �            <, d�            ��( T   �� 
 CResistors��  CValue  � �,     220        �k@      �?   �  x0 �1      t 	        �          �  x@ �A      u 	        �          �  xP �Q      v 	 �v��D/@'�:�?  �  x` �a      w 	        �          �  xp �q      x 	        �          �  x� ��      y 	        �          �  x� ��      z 	        �          �  x� ��      { 	        �          �  �� ��      ^          �          �  �� ��      ]          �          �  �� ��      [          �          �  �p �q      a          �          �  �` �a      b          �          �  �P �Q      c   B��� @'�:��  �  �@ �A      d          �          �  �0 �1      e          �            �, ��            �� v   ��  �� ��     220        �k@      �?   �  x� ��      f          �          �  x� ��      g          �          �  x� ��      h          �          �  x �     i          �          �  x�     j          �          �  x �!     k          �          �  x0�1     l          �          �  x@�A     m          �          �  �@�A     n          �          �  �0�1     o          �          �  � �!     p          �          �  ��     q          �          �  � �     r          �          �  �� ��      s          �          �  �� ��      `          �          �  �� ��      _          �            �� �F     0      �� v   ��  CLED_G�  0 -1      e          �          �  D0 Y1      \                       ,$ DD     B    ��      @��  P -Q      d          �          �  DP YQ      \                       ,D Dd     E    ��      @��  p -q      c   B��� @ �:�?  �  Dp Yq      \            �:��    ,d D�     H  
 ��      @��  � -�      b          �          �  D� Y�      \                       ,� D�     K    ��      @��  � -�      a          �          �  D� Y�      \                       ,� D�     N    ��      @��  P-Q     `          �          �  DPYQ     \                       ,DDd    Q    ��      @��  0-1     _          �          �  D0Y1     \                       ,$DD    T    ��      @��  -     ^          �          �  DY     \                       ,D$    W    ��      @��  � -�      ]          �          �  D� Y�      \                       ,� D    Z    ��      @��  � -�      [          �          �  D� Y�      \                       ,� D�     ]    ��      ��  CSPST��  CToggle  x � 0     `   �  h } 	     Y 	       @          �  � � 	     S         @            | �      c     ��    ��  CBattery�  4 �\ �    5V         @      �? V �  T i 	     Y         @          �  ( = 	     Z                       < �T     h    ��      ��  CClock�  ��     X                       ��    l    ����     �� 
 CCounter10�  01%      S         @          �  %      X                     �  �89     W          �          �  D	Y     )         @          �  DY     R          �          �  (D)Y     Q          �          �  8D9Y     *         @            $<D    o      ��  ,   m��  ��%      S         @          �  `a%      +         @          �  @8U9     W          �          �  XDYY     W          �          �  hDiY     V          �          �  xDyY     U         @          �  �D�Y     T          �            T$�D    w      ��  ,   ��  C4511�  �p��      T          �          �  xpy�      U         @          �  hpi�      V          �          �  XpY�      W          �          �  HpI�      S         @          �  8p9�      S         @          �  (p)�      \                     �  (�)�     2   |��.@�W�/�1��  �  8�9�     1   |��.@�W�/�1��  �  H�I�     0          �          �  X�Y�     /   |��.@�W�/�1��  �  h�i�     .   |��.@�W�/�1��  �  x�y�     -   |��.@�W�/�1��  �  ����     ,          �             ���    �      ��  h   ~��  8x9�      *         @          �  (x)�      Q          �          �  x�      R          �          �  x	�      )         @          �  �x��      S         @          �  �x��      S         @          �  �x��      \                     �  ����     N          �          �  ����     M          �          �  ����     L   {��.@�W�/�1��  �  �	�     K   {��.@�W�/�1��  �  ��     J   {��.@�W�/�1��  �  (�)�     I   {��.@�W�/�1��  �  8�9�     H   {��.@�W�/�1��    ��<�    �      ��  h   ��  ����    220          �k@      �?   �  8�9�      H 	 {��.@�W�/�1�?  �  (�)�      I 	 {��.@�W�/�1�?  �  ��      J 	 {��.@�W�/�1�?  �  �	�      K 	 {��.@�W�/�1�?  �  ����      L 	 {��.@�W�/�1�?  �  ����      M 	        �          �  ����      N 	        �          �  ����      O          �          �  ���     P          �          �  ���     C          �          �  ���     B          �          �  ���     A   �i�n� @�W�/�1��  �  �	     @   �i�n� @�W�/�1��  �  �     G   �i�n� @�W�/�1��  �  (�)     F   �i�n� @�W�/�1��  �  8�9     E   �i�n� @�W�/�1��    ��<�    �      �� v   ��  CSevenSegmentDisplay�  �@�A     @   �i�n� @ W�/�1�?  �  �P�Q     A   �i�n� @ W�/�1�?  �  �`�a     B          �          �  �p�q     C          �          �  |	�     ?           �l��~��  �  $p9q     D          �          �  $`9a     E   �i�n� @ W�/�1�?  �  $P9Q     F   �i�n� @ W�/�1�?  �  $@9A     G   �i�n� @ W�/�1�?    �<$|     � 	     ��0 <            ��  CEarth�  �	�      ? 	         �l��~�?    ���     �    ��      ���  ����     \            �:�?    ����    �    ��      ���  X�Y�      < 	         �l��~�?    K�c�     �    ��      ���  08E9     8   �i�n� @ W�/�1�?  �  0HEI     7          �          �  0XEY     6   �i�n� @ W�/�1�?  �  0hEi     5   �i�n� @ W�/�1�?  �  XtY�     <           �l��~��  �  th�i     =          �          �  tX�Y     ;          �          �  tH�I     :   �i�n� @ W�/�1�?  �  t8�9     9   �i�n� @ W�/�1�?    D4tt     � 	     ��0 <             ��  � ��    220          �k@      �?   �  ����      , 	        �          �  x�y�      - 	 |��.@�W�/�1�?  �  h�i�      . 	 |��.@�W�/�1�?  �  X�Y�      / 	 |��.@�W�/�1�?  �  H�I�      0 	        �          �  8�9�      1 	 |��.@�W�/�1�?  �  (�)�      2 	 |��.@�W�/�1�?  �  ��      3          �          �  ��     4          �          �  (�)�     5   �i�n� @�W�/�1��  �  8�9�     6   �i�n� @�W�/�1��  �  H�I�     7          �          �  X�Y�     8   �i�n� @�W�/�1��  �  h�i�     9   �i�n� @�W�/�1��  �  x�y�     :   �i�n� @�W�/�1��  �  ����     ;          �            ���    �      �� v   ��  CAND�  ��-      )         @          �  ��-      *         @          �  �D�Y     +         @            �,�D    �      ��        �   �     ���  CWire  � ` )a      + �  � ` � 1      + �  � 0Q1     + ��� 
 CCrossOver  N�T�        P0Q�      + �  P�a�     + ��  N�T�      �  ����        @���     W �  ���     \ �   ��      \ �   ���     \ �  �P��      \ �  X�     \ �  � P )Q      S �  � P �       S �  �  �      S ��  �        �  9     S �  �A�     W �  (`)q      \ �  8XIY     S ��  F\Ld        HXIq      S ��  F\Ld      �  �\�d      �  v\|d      �  f\ld      �  V\\d        (`�a     \ ��  V\\d        XXYq      W ��  f\ld        hXiq      V ��  v\|d        xXyq      U ��  �\�d        �X�q      T �  �0 1      e �  �@ A      d �  @ Q       d �  �P Q      c �  p q      c �  P q       c �  �` 	a      b �  � �      b �  ` 	�       b �  �p q      a �   � �      a �   p �       a �  �� ��      [ �  �� ��       [ �  �� �      [ �  �� ��      ] �  �� �      ] �  �� ��       ] �  �� ��      ^ �  �     ^ �  �� ��      _ �  �01     _ �  �� �      ^ �  �� �1      _ �  �� ��      ` �  �� �Q      ` �  �PQ     ` �  X0 �1      \ �  XP �Q      \ �  �0 �Q       \ �  Xp �q      \ �  �P �q       \ �  X� ��      \ �  �p ��       \ �  X� ��      \ �  �� ��       \ �  X� ��      \ �  �� ��       \ �  X� ��      \ �  �� ��       \ �  �� �      \ �  X0�1     \ �  ��1      \ �  XP�Q     \ �  �0�Q      \ �  X� Y�       f �  X� y�      f �  H� I�       g �  H� y�      g �  P�Qa      * ��  6L<T        8 9Y      S �  �  � 	      S ��  �        �Q      W �  PXYY     W �  PPQY      W ��  6L<T        PQQ     W ��  >�D        @�A9      W �       X ��  �      �  ��        �      X ��  �      �  ���      �  ���      �  ���      �  ���        � 1     S ��  ��        ��Q�     * ��  ^�d        `�a      + ��  >�D      �  ^�d        8 �     S �  � �      S �  8`Ya     E �  8 Y     E �  ( )      F �  (Q     F �  X Ya      E �  8PQQ     F �         G �  I     G �  PQQ      F �  HIA      G �  8@IA     G �   	1      @ �  �0	1     @ �  �0�A      @ �  �@�A     @ �  �P�Q     A �  �(�Q      A �  � �)      A �  �`�a     B �  � �a      B �  �(�)     A �  � �!     B �  � �!      B �  �p�q     C �  ��     C �  � �      C ��  dl        X	y      ) ��  dl        Xy      R ��  &d,l        (X)y      Q ��  6d<l      �  &d,l      �  dl      �  dl        �hIi     S �  0 1      S �  0 I     S �  �h�y      S �  �x�y     S �  ��q      C �  (�)      5 �  )     5 �  i      5 �  h1i     5 �  8�9      6 �  9     6 �    I!     7 �  Y      6 �  X1Y     6 �  H�I!      7 �    !I      7 �   H1I     7 �  (819     8 �  (()9      8 �  ((Y)     8 �  X�Y)      8 �  �8�9     9 �  ��9      9 �  ��I      : �  h�     9 �  h�i      9 �  �H�I     : �  ���Y      ; �  x�	     : �  x�y	      : �  ����     ; �  �X�Y     ; �  �`�y      \ �  8pIq     S �  ��Y      ) �  �X	Y     ) ��  ��        ��     ) �  ��      * ��  ���        ���      * ��  F\Ld        H Ii      S ��  F\Ld        8`Qa     * �  8X9a      * ��  6d<l        8`9y      * �  �X�Y     + ��  ���        ���Y      + �  `���     + ��  ����      �  ��      �  ��      �  ���        ���a      \ ��  ��      �  ��        ��     * ��  ��      �  ���        ���9      W     �   �     �    �   �         �   �      �   �        :  8  %   $   #   "   !                      !  ! "  " #  # $  $ %  % & & ' ' ( ( ) ) * * + + , , - - 0 90 1 ;1 2   2 3   3 4   4 5   5 6   6 7   7 8 8   9 9   : :   ; ;   < <   = =   > > #? ? B B C C &E E F F 'H H I I )K K L L +N N O O -Q %Q R R 6T  T U U 4W W X X � Z Z [ [ 1] ] ^ ^ /c h c d d ?h h c i   i l l Io o p Hp q �q r r ts s vt t xu u �w Yw x Tx y Fy z z { { | | } } 	� 	� � � � � � � � �� � �� � � � � � � � � � � � � � � � � � � � � � � � � � �� � x� � v� � t� � �� � �� � �� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �   � � �   � � s� � p� � k� � e� � `� � \� � [� h� � i� � l� � q� � � � � �   � � Z� � _� � d� � � � � �� � � � �� � �� � �� � �� � � � � �   � � �� � �� � �� � � � � � � � � � � � � � � � � � � � � �   � � �   � � �� � �� � �� � �� � �� � �� � �� �� � �� � � ��  � � � � � � � � � �� � � �� �� � � � � � 6� X 5�  � � ?� � A� =@F� � =� � � � � � � � 
� � � � �B� { �  | � 	� } � - B , E + H * K ) N ( ] ' Z & !!W ? ""T  > $#%$Q C (F *&'I ,()L .*+O 0,-^ 2./[ 3012� U 734R 75�  980  ;:1 R�=EV� � d @� � DCz DBD>@CFW� y p IIMISl HLJL�L�L�L�VRK�<TX� x VGVU� YLw � ^� ^� ]\b[Z� b� a`c]_ad� c� fgefhg� j� ni� nm� oljkmp� o�� �s� rt~�� v}s � x|t � z�zyzwzu���o L�z�� � rq� ������� � ��������� � ����� �� ����� �� �������� �� ������ �� �� ��� � � ���r ��� ��� �PR����z���<u ��{�� �� �O��T��� �����Q� � ���������N� q  |          �$s�        @     +        @            @    "V  (      ��                
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 