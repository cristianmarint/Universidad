��  CCircuit��  CSerializeHack           ��  CPart    0   0     ���  CECapacitor��  CValue  ���    100�F(    -C��6?      �?�F �� 	 CTerminal  ��         ���	�I@ɒ)d,`?  �  �                ɒ)d,`�    ��        ��      F�L0ү:?�� 
 CCounter10�  ��	              @          �  �(�)        </��`@          �  �4�I               �          �  �0�1        �o�� @ X�F�Ċ�  �  � �!               �          �  ��               �          �  � �     
          �            �� �4           ��  ,   ��  CLED�  ����       	        �          �  ����                            ����         ��      ��  p�q�       	        �          �  p�q�                            d���         ��      ��  P�Q�       	        �          �  P�Q�                            D�d�          ��      ��  0�1�       	 �g:.��? X�F�Ċ?  �  0�1�                 X�F�Ċ�    $�D�     #  
 ��      �� 
 CResistors
�  	i)w    220          �k@      �?   �  �P�e                �          �  �P�e      
          �          �  �P�e                �          �  pPqe                �          �  `Pae                �          �  PPQe                �          �  @PAe                �          �  0P1e         �o�� @#X�F�Ċ?  �  0|1�        �g:.��?#X�F�Ċ�  �  @|A�               �          �  P|Q�               �          �  `|a�               �          �  p|q�               �          �  �|��               �          �  �|��               �          �  �|��               �            *d�|    (      �� v   �� 	 CPushMake��  CKey  �Z�v      9   �  �t��              @          �  �H�]       	        �            �\�t    <      ��    ��  CBattery
�  !3/    5V(          @      �? V �  @A               @qE�ؑ.��  �  @4AI                qE�ؑ.�?    4L4     A    ��      ��  CEarth�  @HA]       	         qE�ؑ.��    3\Kd     E    ��      ��  CSPST��  CToggle  ��0     G   �  ��	              @qE�ؑ.�?  �  ��	              @qE�ؑ.��    ��     J     ��    �� 	 CResistor
�  ���    220          �k@      �?   �  ��       	 �P��@9 @Aj~�?  �  �                9 @Aj~��    ��     O    ��      ��  CLED_G�  ��         </��`@ !@Aj~�?  �  ��        �P��@ !@Aj~��    �$�     S  
 ��      C��  (=                 �qV|֐�?    <D     V    ��      ��  C555�  �(�=               @=W)�?  �  �(�=               @          �  �@�A     	   ���	�I@          �  �P�Q        ���	�I@          �  �`�a        ���	�I@          �  �d�y                N贁Nk�  �  �d�y        ������
@       �  �  �P�Q        </��`@\@Aj~��    �<�d     Y    ��   (   �� 
 CVResistor��  CSlider   t/�     
�  ���    0k     F]t�1�@        k 
   e �  h}      	 	 ���	�I@˒)d,`?  �  ��        ���	�I@˒)d,`�    |�     f    ��      L�
�  �AO    470          `}@      �?   �  (=               @˒)d,`?  �  Ti     	   ���	�I@˒)d,`�    <T     j    ��          0   0     ���  CWire  � �Q      
 m�  � �     
 m�  pqQ       m�  �q      m�  P QQ       m�  � Q!      m�  001Q       m�  �011      m�  �(�Q       m��� 
 CCrossOver  fLlT        P�Q      m�x�  fLlT        hi�       m�  h�	      m�  Pq      m�  p�      m�  ���       m�  0Q      m�  p�q       m�  1      m�  P�Q       m�  �      m�  0�1       m�          m�  �i	      m�  �	      m�  h���      m�  �      m�  �x�       m�  �	      m�  @�	      m�  )       m�         m�  P�       m�  �PQ      m�  p`q�       m�  pPqa       m�  p`�a      m�  hai     	 m�  ��       m�  ��       m�  �q�      m�  pP�Q      m�  `@ai      	 m�  `@�A     	 m�  ��)       m�  ��	      m�  ��)       m�  )           0   0     �    0   0         0   0      �    �  |   v    =   u   s   q   o  6      4    �   2   ! ! � # 0 # $ $ � (   ( ) n ) *   * + p + ,   , - r - .   . / t / 0 0 # 1 1   2 2   3 3   4 4  5 5   6 6  7 7   < < � =  = A � A B B E E B E J � J K K � O T O P P � S � S T T O V � V Y � Y Z � Z [ � [ \ � \ ] � ] ^ ^ � _ _   ` ` � f k f g g � j � j k k � o )  n q +  p s -  r u /  t  w w { � v z y | � �  � � }   ~ � �  ~ � � ! } � � $ � P � � z � � z < � � ^ � K � A J � V  � w S ` � � � � � � ] f � �  g � � � � \ � � � [ � Y � � � Z � j            �$s�        @     +        @            @    "V  (      �P                
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 