��  CCircuit��  CSerializeHack           ��  CPart    0   0     ���  CECapacitor��  CValue  � ��    100�F(    -C��6?      �?�F �� 	 CTerminal   p!�         �H���?ʒ)d,`�  �   �!�                ʒ)d,`?    �,�        ��      q��gC��>��  CSevenSegmentDisplay�  �� ��                �          �  �� ��                �          �  � �               �          �  ��               �          �  1                @A�c=墿  �  ,A               �          �  , A        �i�n� @ W�/�1�?  �  ,� A�         �i�n� @ W�/�1�?  �  ,� A�         �i�n� @ W�/�1�?    �� ,      	     ��0 <             �� 
 CResistors
�  h� ��     220        �k@      �?   �  X� m�       	 |��.@�W�/�1�?  �  X� m�       	 |��.@�W�/�1�?  �  X� m�       	 |��.@�W�/�1�?  �  X� m�       	        �          �  X� m�       	        �          �  X� m�       	        �          �  X m      	        �          �  Xm               �          �  ��     	          �          �  � �               �          �  �� ��                �          �  �� ��                �          �  �� ��                �          �  �� ��         �i�n� @�W�/�1��  �  �� ��         �i�n� @�W�/�1��  �  �� ��         �i�n� @�W�/�1��    l� �           �� v   ��  C4511�  � %�               @          �  � %�               @          �  � %�               @          �  � %�                �          �  � %�               @          �  � %�               @          �   %               �          �  D Y               �          �  D� Y�                �          �  D� Y�                �          �  D� Y�                �          �  D� Y�         |��.@�W�/�1��  �  D� Y�         |��.@�W�/�1��  �  D� Y�         |��.@�W�/�1��    $� D     /      ��  h   �� 	 CResistor
�  � � �     470          `}@      �?   �   � !�                @<s���?�?  �   � !	        �H���?<s���?��    � $�      @    ��      �� 
 CVResistor��  CSlider  0?<     
�  � !/    0k     F]t�1�@        k 
   F �   !       	 �H���?Ȓ)d,`�  �   4!I        �H���?Ȓ)d,`?    ,4     G    ��      ��  C555�  �� ��                @N贁Nk?  �  �� ��                @          �  �� ��         �H���?��8��J�?  �  �� ��         �H���?          �  � �        �H���?          �  ��                ao9 ?��  �  ��     
   ������
@       �  �  �� 	�                �            �� �     K    ��   (   ��  CEarth�   �!�                 �_D��?    �+�     U    ��      ��  CLED_G�    !5                �          �   L!a               �            44L     X    ��      =�
�  �y�    220          �k@      �?   �   `!u       	        �          �   �!�                            t$�     \    ��      ��  CSPST��  CToggle  � � � �      _   �  � � � �               @z(=e�?  �  � � � �               @z(=e��    � � � �      b     ��    S��  P � Q �        	         z(=e��    C � [      e    ��      ��  CBattery
�   � C �     5V(          @      �? V �  P � Q �                @z(=e��  �  P � Q �                 z(=e�?    D � \ �      i    ��      �� 	 CPushMake��  CKey  �� �      l   �  ��)              @          �  �� ��        	        �            �� �    o      ��    �� 
 CCounter10�  �� ��               @          �  �� ��                �          �  �� ��                �          �  �� ��                �          �  �� ��               @          �  �� ��               @          �  �� ��               @            �� ��      s      ��  ,       0   0     ���  CWire�� 
 CCrossOver  ^� d�       }�  v� |�         X� ��       {�   � Y�       {�  X� YA       {�  X@�A      {�  � �A       {�  �       {�  �� �       {�  �� ��        {�  �� �       {�  �� �9       {�  `8�9      {�}�  ^� d�         `� a9       {�  �� a�       {�  `� y�       {�   �!�       {�   ��      {�  0�       {�  � �      {�  � �       {�  ��      {�  � �      {�  �� �       {�  �� ��       {�  �� ��       {�  �� ��        {�  �� ��       {�  �� ��        {�  �� ��       {�  @ Q      {�  P� Q       {�  �� Q�       {�  H� I�        {�  �� I�       {�  @� I�       {�  @� A�        {�  �� A�       {�   � ��       {�  �� �       {�  �� �       {�  �� �       {�  �� �       {�  � !�       {�   � !�        {�  �� ��        {�  �� ��       {�  �� ��        {�  p� ��       {�  p� q	       {�  �� ��       {�   `�a      {�   H!a       {�   `!q       {�   q	      {�  � �      {�  �� �       {�  � �a       {�   � !!       {�   �!�       {�   �!�       {�  P � � �       {�  � � !�       {�  ���       {�   ���      {�  x(�)      {�  ��!�      {�  x� ��       {�}�  v� |�         x� y)       {�  �� ��            0   0     �    0   0         0   0      �    �  �   �   �   �    �       �   �   �  <   ;   :    9   ! 8 ! " 7 " # 6 # $   $ % %   & & � ' ' � ( ( � ) ) � * * � + + � , , � / � / 0 � 0 1 � 1 2 � 2 3 � 3 4 � 4 5 � 5 6 6 # 7 7 " 8 8 ! 9 9   : :  ; ;  < <  @ � @ A A � G A G H H � K � K L � L M � M N � N O � O P P � Q Q   R R � U � U X � X Y Y \ \ Y \ ] ] � b � b c c � e j e i � i j j e o o � p u p s � s t � t u u p v v � w w � x x � y y � | � | � � � � � | � � � � � � 5 � 4 � � � 3 � � � � � ~ � � � � � � ] � � �  � & � � � �  �  � � ' � �  � � ( � �  ) �  � � � , � � � + �  � �  * � � � v 2 w 1 x 0 y / R � � @ � L � � � K � M � � � N � � H � �  G � � O � � � � � X  � � U i b c � P � � � � o � � � s �  � � t |             �$s�        @     +        @            @    "V  (      �P                
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 