��  CCircuit��  CSerializeHack           ��  CPart�� 
 CTextLabel  )�Q�    Decodi.          �   �     ���  CAND�� 	 CTerminal  �h�}      .          �          �  �h�}      1          �          �  ����     2          �            �|��          ��    �� 
 CResistors��  CValue  )!I/    220          �k@      �?   �  ��      = 	 |��.@�W�/�1�?  �  ��      < 	 |��.@�W�/�1�?  �  ��      ; 	 |��.@�W�/�1�?  �  ��      : 	        �          �  ��      9 	 |��.@�W�/�1�?  �  pq      8 	 |��.@�W�/�1�?  �  `a      7 	 |��.@�W�/�1�?  �  PQ      Y          �          �  P4QI     Z          �          �  `4aI     T   �i�n� @�W�/�1��  �  p4qI     S   �i�n� @�W�/�1��  �  �4�I     R   �i�n� @�W�/�1��  �  �4�I     Q          �          �  �4�I     X   �i�n� @�W�/�1��  �  �4�I     W   �i�n� @�W�/�1��  �  �4�I     V   �i�n� @�W�/�1��    J�4          �� v   ��  CSevenSegmentDisplay�  h�}�     Q          �          �  h�}�     R   �i�n� @ W�/�1�?  �  h�}�     S   �i�n� @ W�/�1�?  �  h�}�     T   �i�n� @ W�/�1�?  �  ����     P           @A�c=岿  �  ����     U          �          �  ����     V   �i�n� @ W�/�1�?  �  ����     W   �i�n� @ W�/�1�?  �  ����     X   �i�n� @ W�/�1�?    |���     & 	     ��0 <           ��  CEarth�  ����      P 	         @A�c=�?    ����     1    ��      /��  �      6                       � �     3    ��      /��  @�A�      N 	          W�/�1�?    3�K�     5    ��      $��  �-�     J   �i�n� @ W�/�1�?  �  �-�     I   �i�n� @ W�/�1�?  �  �-�     H          �          �  �-�     G          �          �  @�A�     N            W�/�1��  �  \�q�     O          �          �  \�q�     M   �i�n� @ W�/�1�?  �  \�q�     L   �i�n� @ W�/�1�?  �  \�q�     K          �            ,�\�     7 	     ��0 <            ��  �)�7    220          �k@      �?   �  pq%      D 	 |��.@�W�/�1�?  �  `a%      C 	 |��.@�W�/�1�?  �  PQ%      B 	        �          �  @A%      A 	 |��.@�W�/�1�?  �  01%      @ 	 |��.@�W�/�1�?  �   !%      ? 	        �          �  %      > 	        �          �   %      E          �          �   <Q     F          �          �  <Q     G          �          �   <!Q     H          �          �  0<1Q     I   �i�n� @�W�/�1��  �  @<AQ     J   �i�n� @�W�/�1��  �  P<QQ     K          �          �  `<aQ     L   �i�n� @�W�/�1��  �  p<qQ     M   �i�n� @�W�/�1��    �$t<    B      �� v   ��  C4511�  p�q�      1          �          �  `�a�      0          �          �  P�Q�      /         @          �  @�A�      .          �          �  0�1�      *         @          �   �!�      *         @          �  ��      6                     �  �     >          �          �   �!     ?          �          �  0�1     @   |��.@�W�/�1��  �  @�A     A   |��.@�W�/�1��  �  P�Q     B          �          �  `�a     C   |��.@�W�/�1��  �  p�q     D   |��.@�W�/�1��    �t�    T      ��  h   R��  ����      5          �          �  ����      4          �          �  ����      3          �          �  ����      -          �          �  ����      *         @          �  p�q�      *         @          �  `�a�      6                     �  `�a	     7   |��.@�W�/�1��  �  p�q	     8   |��.@�W�/�1��  �  ���	     9   |��.@�W�/�1��  �  ���	     :          �          �  ���	     ;   |��.@�W�/�1��  �  ���	     <   |��.@�W�/�1��  �  ���	     =   |��.@�W�/�1��    X���    c      ��  h   �� 
 CCounter10�  �`�u      *         @          �  �`�u      2          �          �  x���     -          �          �  ����     -          �          �  ����     3          �          �  ����     4          �          �  ����     5          �            �t��    s      ��  ,   q��  h`iu      *         @          �  H`Iu      ,                     �  (�=�     -          �          �  @�A�     .          �          �  P�Q�     /         @          �  `�a�     0          �          �  p�q�     1          �            <tt�    {      ��  ,   ��  CClock�  PQ)     ,                       L� T    �    ����     ��  CBattery�  l ?� M    5V         @      �? V �  � X� Y     )         @          �  ` Xu Y     +                       t L� d    �    ��      ��  CSPST��  CToggle  � `� �     �   �  � X� Y     ) 	       @          �  � X� Y     *         @            � T� \     �     ��        �   �     ���  CWire�� 
 CCrossOver  &\,d      ��  &L,T        ()�      - ����  &\,d      ��  \d        �`1a     1 ����        ��  \d      ��  dl      ��  LT         �      6 ��  �0�1     2 ����  �L�T        �0��      2 ��  ����     2 ����  n�t�        p�q�      1 ��  p�q�      1 ����  ~���        p���     1 ����  ~���        �P��      * ����  .L4T        0H1a      1 ��  �`�i      1 ����  dl        �hi     . ��  �A�     . ��  h�      . ��  p���     * ��  ��      6 ��  ����     V ��  �H�I     V ��  �H�Y      W ��  �X�Y     W ��  �H��      V ��  ����     W ��  �H�a      X ��  �`�a     X ��  �X��      W ��  �`��      X ��  ����     X ��  �H�y      Q ��  `x�y     Q ��  `xa�      Q ��  `�i�     Q ��  X�i�     R ��  XpY�      R ��  �H�q      R ��  P�i�     S ��  PhQ�      S ��  Xp�q     R ��  Phqi     S ��  pHqi      S ��  H�i�     T ��  H`I�      T ��  H`aa     T ��  `Haa      T ��  �h��      G ��   �1�     * ��  0�1�      * ��  hP�Q     * ��  hPia      * ����  n�t�      ��  ^�d�      ��  N�T�      ��  >�D�        0���     * ����  ^�d�        `�a�      0 ����  N�T�        P�Q�      / ����  >�D�        @�A�      . ��  Pi      G ��  �hi     G ��  ���     G ��   P!q      H ��   p!q     H ��  x1y     I ��   p�      H ��   ��     H ��  0P1y      I ��  x	�      I ��  ��     I ��  ��     J ��  ��      J ��  �A�     J ��  @PA�      J ��  p���     K ��  �h��      K ��  �`��      L ��  Ph�i     K ��  PPQi      K ��  p���     L ��  �P��      M ��  ``�a     L ��  `Paa      L ��  pP�Q     M ��  p���     M ��  �P�a      * ����  vL|T      ��  �L�T        pP�Q     * ����  �L�T        �0�a      2 ����  NDTL        0H�I     1 ����  NLTT      ��  &L,T      ��  �L�T      ��  .L4T      ��  LT        �PiQ     * ����  NLTT      ��  NDTL        P(Qa      , ��  H`Qa     , ����  n�t�        H���     - ��  ����      - ��  ����     - ��  � P� Y      * ����  n�t�        pPq�      * ��  �H��      1 ����  ����        ����      5 ����  ����        ����      4 ����  ����        ����      3 ����  ����        ����      - ����  ~���      ��  ����      ��  ����      ��  ����      ��  ����        `��     6 ����  ~���        ����      * ��  p���     * ��  `�a�      6 ��  Hy	     - ����  FLLT        � PqQ     * ����          x)	     - ����  vL|T        xy�      - ����  FLLT        HI�      -     �   �     �    �   �         �   �      �   �    �  p   o   n   m   l   k   j            �   �   �     � ! ! � " " � # # � & � & ' � ' ( � ( ) � ) * * 1 + +   , , � - - � . . � 1 * 1 3 3 � 5 ; 5 7 � 7 8 � 8 9 � 9 : � : ; ; 5 < <   = = � > > � ? ? � B a B C ` C D _ D E ^ E F ] F G \ G H [ H I   I J J   K K � L L � M M � N N � O O � P P � Q Q � T � T U � U V � V W � W X � X Y � Y Z � Z [ [ H \ \ G ] ] F ^ ^ E _ _ D ` ` C a a B c c d d e e f f g � g h � h i "i j j  k k  l l  m m  n n  o o  p p  s � s t � t u (u v v w w x x y y { � { | | } � } ~ ~ �   � � � � � � � � � � � � �   � � � � � � � � � &} � � � � � � � '� � � � � 3 � � � � � �  � � � T � � � � � � � � � � � � �  � �  � � ~ � � h � Z , � # � " � � � � � - � ! � � � � � � � . �   � � � � � � & � ' � �  � � ( � � � � � �  � � ) � � � �  � � � Y X � � � � � { � � � � � � � � � � � � � U � �  V � � � W K � � � � : L � � � � � � � � 9 M � � � � 8 � 7 � � � � N � ? � � � � � � � O � > � � � � � P � Q � = � � s � )� � $� � � � t � � � � � � � � � � � � �  � � | 	*	v $� 
� !� � y c x d w e f  "� !g i *($+&� #� (� &u *%#	 [          �$s�        @     +        @            @    "V  (      ��                
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 