��  CCircuit��  CSerializeHack           ��  CPart�� 
 CTextLabel  �� �     CI 555 generador de pulsos          0   0     ���  CECapacitor��  CValue  ���    100�F(    -C��6?      �?�F �� 	 CTerminal  ��         �x�I�Y@�~S%]��>  �  �     
           �~S%]���    ��        ��      �䅻>�/?��  CBattery�  !3/    5V(          @      �? V �  @A               @�g�n�/��  �  @4AI                �g�n�/�?    4L4         ��      ��  CEarth�  @HA]       	         �g�n�/��    3\Kd         ��      ��  CSPST��  CToggle  ��0        �  ��	              @�g�n�/�?  �  ��	              @�g�n�/��    ��          ��    �� 	 CResistor�  ���    220          �k@      �?   �  ��       	 �P��@9 @Aj~�?  �  �     
           9 @Aj~��    ��     "    ��      ��  CLED_G�  ��         </��`@ !@Aj~�?  �  ��        �P��@ !@Aj~��    �$�     &  
 ��      ��  �x��       	         N贁Nk?    ����     )    ��      ��  (=      
           ���o⋉?    <D     +    ��      ��  C555�  �(�=               @=W)�?  �  �(�=               @          �  �@�A     	   -^?���@          �  �P�Q        �x�I�Y@          �  �`�a        �x�I�Y@          �  �d�y                N贁Nk�  �  �d�y        ������
@       �  �  �P�Q        </��`@\@Aj~��    �<�d     .    ��   (   �� 
 CVResistor��  CSlider   t/�     �  ���    100k          j�@      �?k 
   : �  h}      	 	 -^?���@�~S%]��>  �  ��        �x�I�Y@�~S%]���    |�     ;    ��      ��  �AO    470          `}@      �?   �  (=               @uS%]��>  �  Ti     	   -^?���@uS%]���    <T     ?    ��          0   0     ���  CWire  �	      B�  �	      B�  @�	      B�  )      
 B�        
 B�       
 B�         
 B�  P�       B�  �PQ      B�  p`q�       B�  pPqa       B�  p`�a      B�  hai     	 B�  ��       B�  ��       B�  �q�      B�  pP�Q      B�  `@ai      	 B�  `@�A     	 B�  ��)       B�  ��	      B�  ��)       B�  )           0   0     �    0   0         0   0      P    G  E         E    D " ' " # # I & J & ' ' " ) 3 ) + F + . V . / X / 0 U 0 1 S 1 2 N 2 3 3 ) 4 4   5 5 K ; @ ; < < Q ? Y ? @ @ O Y W  C   G +  H F I # H K & 5 J M R S N L 2 ; T Q  < R P L M 1 U O T 0 W . X V C / D ?            �$s�        @     +        @            @    "V  (      �P                
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 