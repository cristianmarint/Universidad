��  CCircuit��  CSerializeHack           ��  CPart�� 
 CTextLabel  1�Y�    Decodi.      �  �� �     CI 555 generador de pulsos          0   0     ���  CECapacitor��  CValue  ���    100�F(    -C��6?      �?�F �� 	 CTerminal  ��         �H���?ʒ)d,`�  �  �     R           ʒ)d,`?    ��        ��      q��gC��>�� 
 CResistors�  �1�    220          �k@      �?   �  ����      d 	 |��.@�W�/�1�?  �  ����      c 	 |��.@�W�/�1�?  �  ����      b 	        �          �  x�y�      a 	        �          �  h�i�      ` 	        �          �  X�Y�      _ 	        �          �  H�I�      ^ 	        �          �  8�9�      Q          �          �  8�9�     N          �          �  H�I�     h          �          �  X�Y�     g          �          �  h�i�     f          �          �  x�y�     e          �          �  ����               �          �  ����     k   �i�n� @�W�/�1��  �  ����     j   �i�n� @�W�/�1��    2���          �� v   ��  CSevenSegmentDisplay�  P e!     e          �          �  P0e1     f          �          �  P@eA     g          �          �  PPeQ     h          �          �  x\yq     V            W�/�1��  �  �P�Q     i          �          �  �@�A     j   �i�n� @ W�/�1�?  �  �0�1     k   �i�n� @ W�/�1�?  �  � �!               �            d�\     ' 	     ��0 <             ��  C4511�  �X�m      \         @          �  �X�m      [          �          �  �X�m      Z          �          �  xXym      Y          �          �  hXim      W         @          �  XXYm      W         @          �  HXIm      R                     �  H�I�     ^          �          �  X�Y�     _          �          �  h�i�     `          �          �  x�y�     a          �          �  ����     b          �          �  ����     c   |��.@�W�/�1��  �  ����     d   |��.@�W�/�1��    @l��    2      ��  h   �� 
 CCounter10�  ���      W         @          �  ���      U 	        �          �  ` u!     $          �          �  x,yA     Y          �          �  �,�A     Z          �          �  �,�A     [          �          �  �,�A     \         @            t�,    B      ��  ,   ��  CEarth�  xpy�      V 	          W�/�1�?    k���     K    ��      ��  CAND�  ����      S          �          �  x�y�      T          �          �  ����     U          �            t���    N      ��    L��  �0�E               @          �  �0�E                �          �  �\�q     
          �            �D�\    R      ��    I��  ����      L 	         @A�c=�?    ���     V    ��      @��  �p��      W         @          �  �p��      
 	        �          �  ����     $          �          �  ����     S          �          �  ����     P          �          �  ����     O          �          �  ����     T          �            ����    X      ��  ,   0��  ����      T          �          �  ����      O          �          �  ����      P          �          �  ����      S          �          �  ����      W         @          �  ����      W         @          �  ����      R                     �  ��     B   |��.@�W�/�1��  �  ��     A   |��.@�W�/�1��  �  ��     @   |��.@�W�/�1��  �  ��     ?          �          �  ��     >   |��.@�W�/�1��  �  ��     =   |��.@�W�/�1��  �  ��     <   |��.@�W�/�1��    ���    `      ��  h   %��  ����     H          �          �  ����     G   �i�n� @ W�/�1�?  �  ����     F   �i�n� @ W�/�1�?  �  ����     E   �i�n� @ W�/�1�?  �  ����     L           @A�c=岿  �  ����     M          �          �  ����     K   �i�n� @ W�/�1�?  �  ����     J   �i�n� @ W�/�1�?  �  ����     I   �i�n� @ W�/�1�?    ����     o 	     ��0 <           ��  Y1y?    220          �k@      �?   �  ��-      < 	 |��.@�W�/�1�?  �  ��-      = 	 |��.@�W�/�1�?  �  ��-      > 	 |��.@�W�/�1�?  �  ��-      ? 	        �          �  ��-      @ 	 |��.@�W�/�1�?  �  ��-      A 	 |��.@�W�/�1�?  �  ��-      B 	 |��.@�W�/�1�?  �  ��-      C          �          �  �D�Y     D          �          �  �D�Y     E   �i�n� @�W�/�1��  �  �D�Y     F   �i�n� @�W�/�1��  �  �D�Y     G   �i�n� @�W�/�1��  �  �D�Y     H          �          �  �D�Y     I   �i�n� @�W�/�1��  �  �D�Y     J   �i�n� @�W�/�1��  �  �D�Y     K   �i�n� @�W�/�1��    z,�D    z      �� v   �� 	 CPushMake��  CKey  H� l�       �   �  8� M�      W         @          �  d� y�      $          �            L� d�      �      ��    L��    5               @          �  � �5               @          �  �L�a              @            �4L    �      ��    ��  1�Q�    220          �k@      �?   �  ����      " 	 |��.@�W�/�1�?  �  ����      4 	 {��.@�W�/�1�?  �  ����       	 |��.@�W�/�1�?  �  ����       	 |��.@�W�/�1�?  �  ����       	        �          �  x�y�       	        �          �  h�i�      . 	 |��.@�W�/�1�?  �  X�Y�                �          �  X�Y               �          �  h�i     9   �i�n� @�W�/�1��  �  x�y     8          �          �  ���     7          �          �  ���     6   �i�n� @�W�/�1��  �  ���     !   �i�n� @�W�/�1��  �  ���        �i�n� @�W�/�1��  �  ���     ;   �i�n� @�W�/�1��    R���    �      �� v   %��  p@�A     6   �i�n� @ W�/�1�?  �  pP�Q     7          �          �  p`�a     8          �          �  pp�q     9   �i�n� @ W�/�1�?  �  �|��     5           �l��~��  �  �p�q     :          �          �  �`�a     ;   �i�n� @ W�/�1�?  �  �P�Q        �i�n� @ W�/�1�?  �  �@�A     !   �i�n� @ W�/�1�?    �<�|     � 	     ��0 <             I��  ����      5 	         �l��~�?    ����     �    ��      I��  � �                              � $�     �    ��      I��  H�I�      3 	         �l��~�?    ;�S�     �    ��      %��   H5I     /   �i�n� @ W�/�1�?  �   X5Y        �i�n� @ W�/�1�?  �   h5i               �          �   x5y     %          �          �  H�I�     3           �l��~��  �  dxyy     &          �          �  dhyi     2   �i�n� @ W�/�1�?  �  dXyY     1   �i�n� @ W�/�1�?  �  dHyI     0   �i�n� @ W�/�1�?    4Dd�     � 	     ��0 <            ��  ���    220          �k@      �?   �  x�y�      ' 	 |��.@�W�/�1�?  �  h�i�      ( 	 |��.@�W�/�1�?  �  X�Y�      ) 	 |��.@�W�/�1�?  �  H�I�      * 	 |��.@�W�/�1�?  �  8�9�      + 	 {��.@�W�/�1�?  �  (�)�      , 	        �          �  ��      - 	        �          �  �	�                �          �  �		               �          �  �	     %          �          �  (�)	               �          �  8�9	        �i�n� @�W�/�1��  �  H�I	     /   �i�n� @�W�/�1��  �  X�Y	     0   �i�n� @�W�/�1��  �  h�i	     1   �i�n� @�W�/�1��  �  x�y	     2   �i�n� @�W�/�1��    �|�    �      �� v   0��  x�y�               @          �  h�i�                �          �  X�Y�                �          �  H�I�               @          �  8�9�      W         @          �  (�)�      W         @          �  ��                            �  ��     -          �          �  (�)�     ,          �          �  8�9�     +   {��.@�W�/�1��  �  H�I�     *   |��.@�W�/�1��  �  X�Y�     )   |��.@�W�/�1��  �  h�i�     (   |��.@�W�/�1��  �  x�y�     '   |��.@�W�/�1��    �|�    �      ��  h   0��  �x��               @          �  �x��               @          �  �x��                �          �  �x��                �          �  �x��      W         @          �  xxy�      W         @          �  hxi�                            �  h�i�     .   |��.@�W�/�1��  �  x�y�               �          �  ����               �          �  ����        |��.@�W�/�1��  �  ����        |��.@�W�/�1��  �  ����     4   {��.@�W�/�1��  �  ����     "   |��.@�W�/�1��    `���    �      ��  h   @��  ��-      W         @          �  ��-               @          �  �@�A     $          �          �  �L�a               �          �  �L�a               �          �  �L�a              @          �  �L�a              @            �,�L    �      ��  ,   @��  pq-      W         @          �  PQ-                �          �  0@EA     $          �          �  HLIa              @          �  XLYa               �          �  hLia               �          �  xLya              @            D,|L    �      ��  ,   ��  CBattery�  !3/    5V(          @      �? V �  @A               @z(=e��  �  @4AI                z(=e�?    4L4        ��      I��  @HA]       	         z(=e��    3\Kd        ��      ��  CSPST��  CToggle  ��0       �  ��	              @z(=e�?  �  ��	     W         @z(=e��    ��         ��    �� 	 CResistor�  ���    220          �k@      �?   �  ��       	        �          �  �     R                       ��        ��      ��  CLED_G�  ��                �          �  ��               �            �$�        ��      I��  �x��       	         ao9 ?�?    ����        ��      I��  (=      R           ʒ)d,`�    <D        ��      ��  C555�  �(�=      W         @N贁Nk?  �  �(�=      W         @          �  �@�A     	   �H���?��8��J�?  �  �P�Q        �H���?          �  �`�a        �H���?          �  �d�y                ao9 ?��  �  �d�y        ������
@       �  �  �P�Q               �            �<�d        ��   (   �� 
 CVResistor��  CSlider   t/�     �  ���    0k     �����F�@        k 
   (�  h}      	 	 �H���?Ȓ)d,`�  �  ��        �H���?Ȓ)d,`?    |�     )   ��      ��  �AO    470          `}@      �?   �  (=      W         @<s���?�?  �  Ti     	   �H���?<s���?��    <T     -   ��          0   0     ���  CWire�� 
 CCrossOver  F<LD        @iA     W 0�  � @A     W 0�  @I      W 0�2�  FDLL      2�  fDlL      2�  vD|L      2�  �D�L      2�  �D�L      2�  �D�L        H�I     W 0�  ���I      W 0�2�  FDLL      2�  F<LD        H(IY      R 0�  ����     W 0�  ��	     W 0�2�  ��        ��	     W 0�2�  �� ��         �� �	      W 0�  � � ��      W 0�2�  �� ��         0� ��      $ 0�  � � � A      W 0�2�  fDlL        h@iY      W 0�  XXiY     W 0�  H()     R 0�  )      R 0�  A     R 0�        R 0�  `�a!      $ 0�2�  >�D�        `���     $ 0�2�  >�D�      2�  >�D�        @A�      R 0�  ���     T 0�2�  ��      2�  ��        �!      T 0�  0 !     T 0�   ���     $ 0�2�  .�4�        0�1!      T 0�2�  .�4�      2�  ����      2�  >�D�        ����     S 0�  x�1�     T 0�  x�y�      T 0�2�  ����        ����      $ 0�  �@�A     j 0�  ����     j 0�  ����      k 0�  ����     k 0�  ���A      j 0�  �0�1     k 0�  ����       0�  ����      0�  ���1      k 0�  ���!       0�  � �!      0�  x�y      e 0�  Hy     e 0�  HI!      e 0�  H Q!     e 0�  @0Q1     f 0�  @A1      f 0�  h�i	      f 0�  8@QA     g 0�  8 9A      g 0�  @i	     f 0�  8 Y     g 0�  X�Y      g 0�  0PQQ     h 0�  0�1Q      h 0�  0�I�     h 0�  H�I�      h 0�2�  vD|L        x@yY      Y 0�2�  �D�L        �@�Y      Z 0�2�  �D�L        �@�Y      [ 0�2�  �D�L        �@�Y      \ 0�  �(�1       0�  �())      0�  (X))       0�2�  vT|\        (X�Y      0�2�  vT|\      2�  v|        xya      W 0�  �X�a       0�  �`�a      0�2�  �d�l      2�  �d�l      2�  �d�l      2�  �d�l      2�  �d�l      2�  �d�l        hhi       0�  x`�a     W 0�  �0I1      0�  H0I�       0�  PQq      9 0�  X Ya      8 0�  H���      0�  �`��       0�  �`�a      0�  �`�a     ; 0�  ���a       0�  ����      0�  � �a      ; 0�2�  �d�l        �`��       0�  � �     ; 0�  ��      0�  ��A      ! 0�  ��     ! 0�  �`�a      0�  �`�a      0�2�  ��      2�  ����      2�  ����      2�  ����      2�  ����        ��9�     W 0�  �p9q     W 0�  @     R 0�  �q�      0�  8�9�      W 0�  8p9�      W 0�2�  ����      2�  ����        ����      T 0�2�  ����      2�  ����        ����      O 0�2�  ����      2�  ����        ����      P 0�2�  ����      2�  ����        ����      S 0�2�  ����        ����      W 0�2�  ��      2�  ����      2�  ����      2�  ����      2�  ����      2�  ����        ��!�     $ 0�   �!�      $ 0�2�  .4      2�  .4      2�  .4        0� 1A      $ 0�  �� ��      $ 0�2�  � �       2�        2�  $      2�        2�          � i        0�  ����     W 0�  `(aQ      7 0�  h0iA      6 0�2�  ~�      2�  .4      2�  ��      2�  ��      2�  6<      2�  v|      2�        2�  ��        Q      0�  @���     R 0�  hhiy        0�  xx�y     W 0�2�  �d�l        �`�y      W 0�2�  �d�l        �`�y       0�  ��Q       0�  ���      W 0�2�  �d�l        ��q      W 0�2�  ��        � �i       0�  8���     W 0�  �X�q      E 0�  xp�q     E 0�  xpy�      E 0�  x���     E 0�  �X�y      F 0�  �x�y     F 0�  ����     G 0�  �x��      F 0�  ����     F 0�  �X��      G 0�  ����      G 0�  ����     G 0�  ����     H 0�  ����      H 0�  ����     H 0�  �X��      H 0�  ���     I 0�   p�      I 0�  h	�      J 0�  �pq     I 0�  �X�q      I 0�  ��	�     J 0�  X�      K 0�  �h	i     J 0�  �X�i      J 0�  �XY     K 0�  ���     K 0�2�  ~�      2�  ~�        �� �A      $ 0�  x� ��      $ 0�2�  ~�      2�  ��        x�	     W 0�2�  � �         �� 1�      $ 0�2�  .4      2�          �9      0�2�  .4      2�  ��      2�  6<      2�          �q	     W 0�  8 �      0�   � 9�      W 0�   � !	      W 0�  �!	     W 0�   y	     W 0�2�  ��      2�  ��        �� �       0�  �� ��       0�2�  ��      2�  ��        �� �a       0�2�  vl|t        xhy�       0�  x`yi       0�2�  �d�l        xh�i      0�2�  6<      2�  6<        8 9       0�  ��!       0�2�  $          !!      0�   `Ia      0�    !a       0�  h�        0�2�  �d�l        �`�y       0�2�  �d�l        �`�y       0�2�  �d�l        �`�y       0�  � �       0�  �P�Q      0�  � �      ! 0�  �@�A     ! 0�  � �1      6 0�  h0�1     6 0�  h@qA     6 0�  `PqQ     7 0�  � �)      7 0�  X`qa     8 0�  `(�)     7 0�  X y!     8 0�  x y!      8 0�  Ppqq     9 0�  Pi     9 0�  h i      9 0�    y      % 0�  p`�a      0�  (�9�     W 0�  8p9�      W 0�  p�	     W 0�  pq      W 0�2�  vl|t      2�  fllt      2�  Vl\t      2�  FlLt        8p�q     W 0�2�  fllt        h`i�       0�2�  Vl\t        X`Y�       0�2�  FlLt        H`I�       0�  !      % 0�    !     % 0�   x!y     % 0�  ())       0�  ())      0�  091      0�  (	i       0�  h!i      0�  891       0�  0Y       0�  X!Y      0�  H!I     / 0�  8I      / 0�  8I9     / 0�  HI9      / 0�  xH�I     0 0�  � �I      0 0�  ��Y      1 0�  X �!     0 0�  XY!      0 0�  xX�Y     1 0�  ��i      2 0�  h�     1 0�  hi      1 0�  x�	     2 0�  xh�i     2 0�  @�	      0�  �	     W 0�  PQ       0�  Q       0�2�  ��        ��      W 0�  �	     W 0�         R 0�  P�       0�  �PQ      0�  p`q�       0�  pPqa       0�  hai     	 0�  ��       0�  ��       0�  pP�Q      0�  `@ai      	 0�  `@�A     	 0�  ��)      W 0�  ��	     W 0�  ��)      W 0�  )      W     0   0     �    0   0         0   0      �   Q ?   >   =   <   ;   :   9            �  ~    y! ! s" " n# # j$ $ i' v' ( w( ) z) * * + + K , ,   - - h. . m/ / r2 �2 3 �3 4 �4 5 �5 6 M6 7 M7 8 >8 9 9  : :  ; ;  < <  = =  > >  ? ?  B AB C P C D RD E E �F F �G G �H H �K + K N `N O eO P P C R �R S �S T T Y V s V X �X Y T Y Z fZ [ [ �\ \ �] ] �^ ^ �` �` a �a b �b c �c d �d e �e f �f g g � h h  i i ~ j j } k k | l l { m m z o o p p q �q r �r s s V t t   u u v v w w z m z { l { | k | } j } ~ i ~  h  � g � �   � � �   � � �� � �� � �� � � � 
� � � � � #� � � � 7� � 6� � � �� � � � � � � � � � � � � � � � � � � � � �   � � �   � � Q� � N� � J� � F� � D� � B� � �� H� � I� � K� � O� � � � � �   � � �� � C� � E� � � � � �� � � � n� � m� � j� � e� � � � � �   � � |� � w� � r� � � � � � � � � � � � � � � � � � � � � �   � � �   � � c� � f� � k� � q� � v� � z� � {� .� � ]� � _� � a� � U� � T� � ;� � � � � � � � � � � � � � � � � � � � � � � <� � >� � @� � �� � �� � �� � �� � � � � � � � � � � � � � � � � � � � � � � �� � '� � � � � �� � @� � >� � <� W� � � � �� � � a� � _� � ]� � 0}}~��!O���� S !!""  ##�).)**�-�-..�1@4KJ5166?6L6�6�6�6�5=A6>7>3N8 B =C�C��EEIGBJEHF��G4K816 7 K>QNOU PSD SVRZ UTUc��^ YY�Y�X\^Y��^ad\`_`g`WN [ e^dO fbS�- l$ l# kjpih. p" onqkmor/ q! tustvu' x( |w  |{) }zxy{~ }�* ��� ��9E 5 �:F 4 �;G 3 �<H 2 �S ����������������� �����=�?�A���;��R ���POMK������� ������������ �B��ED�� �+� �Z����������X �P�����������X` ����] a ����\ b ����`c ���d �[����������f��]����� H]���8���!� �e �LIGH����(�-�5�������Uf �� � ����� ���� �CB��2VX�D"1��� ������r � ��� ����q � �� p o � w 	
� 	v � � u �� � )&��H��63�,4�W3�$� #&�$%�'�'*� '+++�*�.Y0� � 11�.�3 3�"� 7�� ::� 79�� <��� >�� � @�� � � �� �� �� �� G�F�� �� � L�� �J�N� M�� �Q� Pde� � � XTCV� X/X^X`XbU�]Z� � _[� � a\9� � dRcR� � giflkgji� � hhml� o� pnoq� p� surywvs� u� t{|zt� y� x� x��� ����� ����#����S)�� *�������%�~- l          �$s�        @     +        @            @    "V  (      �                
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 