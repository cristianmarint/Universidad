��  CCircuit��  CSerializeHack           ��  CPart�� 
 CTextLabel  �i�w    Pulsos          x   x     ���  CECapacitor��  CValue  �1?    100�F(    -C��6?      �?�F �� 	 CTerminal  -         �JS<���?�9
E�0�  �  DY     
           �9
E�0?    ,D        ��      ˛)��!?�� 	 CPushMake��  CKey  `x��         �  Ppeq              @          �  |p�q               �            dh|t           ��    ��  CEarth�  � �� �      C 	          L�Ir�?    � �� �         ��      �� 
 CResistors�  ��$    220        �k@      �?   �  �(�)     2 	 |��.@�W�/�1�?  �  �8�9     3 	 |��.@�W�/�1�?  �  �H�I     4 	 |��.@�W�/�1�?  �  �X�Y     5 	 |��.@�W�/�1�?  �  �h�i     6 	 |��.@�W�/�1�?  �  �x�y     7 	 |��.@�W�/�1�?  �  ����     8 	 |��.@�W�/�1�?  �  ����     9          �          �  ���     :          �          �  ���     ;   �i�n� @�W�/�1��  �  �xy     <   �i�n� @�W�/�1��  �  �hi     =   �i�n� @�W�/�1��  �  �XY     >   �i�n� @�W�/�1��  �  �HI     ?   �i�n� @�W�/�1��  �  �89     @   �i�n� @�W�/�1��  �  �()     A   �i�n� @�W�/�1��    �$��           �� v   ��  C4511�  x(�)        �v��D/@          �  x8�9               �          �  xH�I               �          �  xX�Y     &   �v��D/@          �  xh�i               �          �  xx�y               �          �  x���     C                     �  ����     8   |��.@�W�/�1��  �  �x�y     7   |��.@�W�/�1��  �  �h�i     6   |��.@�W�/�1��  �  �X�Y     5   |��.@�W�/�1��  �  �H�I     4   |��.@�W�/�1��  �  �8�9     3   |��.@�W�/�1��  �  �(�)     2   |��.@�W�/�1��    �$��     /      ��  h   ��  CSevenSegmentDisplay�  � 8� 9     >   �i�n� @ W�/�1�?  �  � H� I     =   �i�n� @ W�/�1�?  �  � X� Y     <   �i�n� @ W�/�1�?  �  � h� i     ;   �i�n� @ W�/�1�?  �  � t� �     C            L�Ir��  �  � h	i     B          �          �  � X	Y     A   �i�n� @ W�/�1�?  �  � H	I     @   �i�n� @ W�/�1�?  �  � 8	9     ?   �i�n� @ W�/�1�?    � 4� t     ? 	     ��0 <           ��  �x��      /            X�F�Ċ?    ����     I    ��      ��  CLED�  X	m      1 	        �          �  �	�     /                       �l�     L    ��      �� 	 CResistor�  �1?    220          �k@      �?   �  	-      $          �          �  D	Y     1          �            ,D     Q    ��      N��  �1�?    220          �k@      �?   �  ��-      %   �o�� @#X�F�Ċ?  �  �D�Y     0   �g:.��?#X�F�Ċ�    �,�D     U    ��      J��  �X�m      0 	 �g:.��? X�F�Ċ?  �  ����     /            X�F�Ċ�    �l��     X  
 ��      J��  (X)m      '          �          �  (�)�     /                       l<�     [    ��      J��  XXYm      #          �          �  X�Y�     /                       Lll�     ^    ��      J��  �X�m      "          �          �  ����     /                       |l��     a    ��      J��  pXqm                �          �  p�q�     /                       dl��     d    ��      J��  @XAm                �          �  @�A�     /                       4lT�     g    ��      J��  Xm                �          �  ��     /                       l$�     j    ��      J��  �X�m                 �          �  ����     /                       �l��     m    ��      J��  �X�m      !          �          �  ����     /                       �l��     p    ��      ��  �>�L    220        �k@      �?   �  xP�Q               �          �  x`�a               �          �  xp�q               �          �  x���                �          �  x���     !          �          �  x���     "          �          �  x���     #          �          �  x���     '          �          �  ����     (          �          �  ����     )          �          �  ����     *          �          �  ����     +          �          �  ����     .          �          �  �p�q     -          �          �  �`�a     ,          �          �  �P�Q               �            �L��     t      �� v   ��  CDecoder�  p���        �v��D/@          �  p���               �          �  p���               �          �  p���     &   �v��D/@          �  ���	     %   �o�� @ X�F�Ċ�  �  ���	     $          �          �  ����     (          �          �  ����     )          �          �  ����     *          �          �  ����     +          �          �  ����     .          �          �  ����     -          �          �  ����     ,          �          �  ����               �            �|��     �      ��  T   ��  ����                 !�:�?    ����     �    ��      ��  CLED_G�           �v��D/@��:�?  �  4I        �+�う@��:��    $4     �  
 ��      J��  ��                �          �  �4�I               �            �4     �    ��      ��  CLED_Y�  ��                �          �  �4�I               �            ��4     �    ��      ��  �a�o    220          �k@      �?   �   H!]                �          �  H]       	 �+�う@�:�?  �   H]                �          �  �H�]       	        �          �  �H�]                �          �  �H�]       	        �          �  �H�]                �          �  �H�]       	 �+�う@(�:�?  �  �t��                (�:��  �  �t��                          �  �t��                          �  �t��               �          �  �t��                          �   t�               �          �  t�                �:��  �   t!�               �            �\$t    �      �� v   ���  ��      &   �v��D/@��:�?  �  �4�I        �+�う@��:��    ��4     �  
 ��      �� 
 CCounter10�  ����              @          �  ����               �          �  ����               �          �  ���     &   �v��D/@@�:��  �  ���               �          �  ���               �          �  �xy        �v��D/@��:��    �t��     �      ��  ,   N��  93G    220          �k@      �?   �  8 95       	        �          �  8L9a     
                       44<L     �    ��      ���  8�9�                �          �  89!               �            ,�L     �    ��      ��  �p��                 m?��̪�?    ����     �    ��      ��  p�      
           �9
E�0�    ��     �    ��      ��  C555�  �p��               @N贁Nk?  �  �p��               @          �  ����     	   ��WY�L�?�8yG,ׅ?  �  ����        �JS<���?          �  ����        �JS<���?          �  ����                m?��̪��  �  ����        ������
@       �  �  ����               �            ����     �    ��   (   �� 
 CVResistor��  CSlider   �/�     �  ���    5k          j�@�������?k 
   � �  ��      	 	 ��WY�L�?�9
E�0�  �  ��        �JS<���?�9
E�0?    ��     �    ��      N��  ���    470          `}@      �?   �  p�               @��(�R�?  �  ��     	   ��WY�L�?��(�R��    ��     �    ��      ��  CSPST��  CToggle  `���     �   �  P�e�              @�c�2&�?  �  |���              @�c�2&��    d�|�     �     ��    ��  � � %       	         �c�2&��    � $� ,     �    ��      ��  CBattery�  � �� �    5V(          @      �? V �  � �� �               @�c�2&��  �  � ��                 �c�2&�?    � �� �     �    ��          x   x     ���  CWire  �p�q      ��� 
 CCrossOver  ����        �p��       �  ����      ���  ����        X���      �  HpQq      �  HPIq       �  �PIQ      �  HP�Q      �  X�Y�       �  8�9�       �  xXya      & ���  f\ld        X`ya     & ���  f\ld      ��  f�l�      ��  f�l�      ��  fdll        hHi�       ���  V�\�      ��  V�\�        X`Y�      & �  X�Q�     & ���  V�\�      ��  f�l�      ��  ^�d�        � �y�     C ���  V�\�        p �i�      �  P�Q�      & �  P�a�     & �  H�I�       �  @�A�      ; �  8�9y      < �  `�a�      & ���  �$�      ��  &�,�      ��  6�<�      ��  F�L�        `�Y�     & �  X�Y�      & ���  F�L�      ��  6�<�      ��  &�,�         �Y�     & ���  �$�         �!�      & ���  &�,�      ��  &�,�        (�)�       ���  6�<�      ��  6�<�      ��  6�<�        8�9       ���  F�L�      ��  F�L�      ��  F�L�      ��  F�L�        HxI	       �  I	      �  X�q�     & �  P�q�      ���  F�L�      ��  6�<�        (�Q�      ���  N�T�      ��  NtT|      ��  NT$      ��  NT        PQ�       ���  N�T�      ��  F�L�        8�Y�      ���  NtT|      ��  Vt\|      ��  ^td|        Hxqy      ���  NT$      ��  V\$        �  a!      ���  NT        � Y      �  p Q      �  p q �       ���  f�l�        `�I�      ���  ^�d�        `ha�       ���  fdll        `hqi      �  hHyI      �  phqy       �  `aY      A �  HYI     @ �  XYI      @ ���  f�l�      ��  f�l�      ��  f�l�      ��  f�l�      ��  f�l      ��  fl      ��  fl        h�i9       �  X�q�      ���  Vt\|      ��  V\$        XY�       �  � � �       �  � �i�      �  � �y�      �  �  � �       ���  v�|�      ��  v�|�      ��  v�|�      ��  v�|�      ��  v�|      ��  v|      ��  v|        x�y)       ���  f�l�      ��  v�|�        x �A�     ; ���  f�l�      ��  v�|�        � �9�     < ���  f�l�      ��  v�|�        � �1�     = ���  f�l�      ��  v�|�        � �)�     > ���  f�l      ��  v�|        P !     ? ���  fl      ��  v|        `     A �  h8y9      �  `�q�      ���  ^td|        ` a�       ���  fl      ��  v|        X	     @ �  8`9�      
 �  H`I�      
 �  pxyy      �  phyi      �  H�Y�      �  8�Y�      �  � `� i      ; �  x `� a     ; �  x �y a      ; �   �A�     ; �  � P� Y      < �  � P� Q     < �  � �� Q      < �   x9y     < �  � H� I     = �  � �� I      = �  � �� 9      > �  0�1i      = �  (�)Y      > �   h1i     = �  � 8� 9     > �   X)Y     > �  8Q9     ? �  P Q9      ? �    !I      ? �  9      @ �   H!I     ? �  )      A �   89     @ �  XaY     A �   ()     A �  �x�y     / �  �x��      / �  ����     / �  ��	�     / �  �)�     / �  (�Y�     / �  X���     / �  ����     / �  ����     / �  ���     / �  �A�     / �  @�q�     / �  ��      % �  �		     % �  �		      % �       $ �  ��     % �  ��      % �  �      $ �  �)�     % �  ��       �  (�)�      % �  0�1�      $ �  (�1�     % �  0h1�      % ���  6d<l        0hIi     % ���  FTL\        H0Ii      % ���  6d<l        8X9�      $ ���  FTL\        8XYY     $ �  H0�1     % �  ��1      % �  X8�9     $ �  ((!)     ' �  X0)1     # �  �!�     $ �   �!�      $ �   �!)      ' �   �1�     $ �  0�9�     $ ���  6�<�      ��  6�<�      ��  6�<�        8�9A      ! ���  >�D�      ��  >�D�      ��  >�D�      ��  >�D�        @�AI        �  X8YY      $ �  ��9      $ �  (()Y      ' ���  &�,�      ��  .�4�      ��  6�<�      ��  >�D�      ��  F�L�      ��  V�\�      ��  f�l�         �y�     ' ���  &�,�        (�)1      # ���  .�4�      ��  .�4�        0�19      " ���  F�L�      ��  F�L�      ��  F�L�      ��  F�L�      ��  F|L�        HpIQ       ���  V�\�      ��  V�\�      ��  V�\�      ��  V�\�      ��  V|\�      ��  Vl\t        X`YY       ���  f�l�      ��  f�l�      ��  f�l�      ��  f�l�      ��  f|l�      ��  fllt      ��  f\ld        hPiY       �  X0YY      # �  �819     " ���  .�4�      ��  6�<�      ��  >�D�      ��  F�L�      ��  V�\�      ��  f�l�        (�y�     # �  �8�Y      " �  �@9A     ! ���  6�<�      ��  >�D�      ��  F�L�      ��  V�\�      ��  f�l�        0�y�     " �  �@�Y      ! �  �HAI       ���  >�D�      ��  F�L�      ��  V�\�      ��  f�l�        8�y�     ! �  �H�Y        �  PIQ      ���  F|L�      ��  V|\�      ��  f|l�        @�y�       �  PY       �  @XYY      ���  Vl\t      ��  fllt        Hpyq      ���  f\ld        X`ya      �  hXqY      �  hPyQ      �  H�9�     
 �  � �Q�      �  ��1�     ( ���  .�4�      ��  .�4�      ��  .�4�      ��  .|4�      ��  .l4t      ��  .\4d      ��  .L4T        0�1�      ( ���  .�4�        ��9�     ) ���  .�4�      ��  6�<�        ��A�     * ���  .�4�      ��  6�<�      ��  >�D�        ��I�     + ���  .|4�      ��  6|<�      ��  >|D�      ��  F|L�        ��Q�     . ���  .l4t      ��  6l<t      ��  >lDt      ��  FlLt      ��  NlTt        �pYq     - ���  .\4d      ��  6\<d      ��  >\Dd      ��  F\Ld      ��  N\Td      ��  V\\d        �`aa     , ���  .L4T      ��  6L<T      ��  >LDT      ��  FLLT      ��  NLTT      ��  VL\T      ��  ^LdT        �PiQ      �  ��1�     ( ���  6�<�      ��  6�<�      ��  6|<�      ��  6l<t      ��  6\<d      ��  6L<T        8�9�      ) �  ��9�     ) ���  >�D�      ��  >|D�      ��  >lDt      ��  >\Dd      ��  >LDT        @�A�      * �  ��A�     * ���  F|L�      ��  FlLt      ��  F\Ld      ��  FLLT        H�I�      + �  ��I�     + ���  NlTt      ��  N\Td      ��  NLTT        P�Q�      . �  ��Q�     . ���  V\\d      ��  VL\T        X�Yq      - �  ��Y�     - ���  ^LdT        `�aa      , �  ��a�     , �  h�iQ       �  ��i�      �   �!�      & �  (�)�       �  8�9�       �  pxq�       �  xIy      �  ���	      & �  ��!�     & �  ��)�      �  �!�     & �  ���	       �  � 9      �  �)�      �  � �	       �  �9�      �  ����      �  ���      �  ����       �  ����       �  ����      �  ����      �  ����       �  ����      �  ����       �  ����       �  ����       �  q	      �  ���q       �  p���      �  P�Q      �  8�9�       �  �P��       �  p�q	       �  p�q�       �  `q      
 �  Xa      
 �  `Ia     
 �  �a�     	 �  �PQ      �  ��9�      �  �p�q      �         �  �	       �  p���      �  `�a�      	 �  `���     	 �  �P�q       �  �P�Q      �  �P�q       �  Pq       �  �P��       �  ����      �  � �� �           x   x     �    x   x         x   x      �   � �    �  C   <   ;   :    9   ! 8 ! " 7 " # 6 # $   $ % %   & & �' ' �( ( �) ) �* * �+ + �, , �/ _/ 0 y0 1 J1 2 � 2 3 �3 4 �4 5 5 6 6 # 7 7 " 8 8 ! 9 9   : :  ; ;  < <  ? �? @ �@ A �A B �B C C D D   E E �F F MG G �I �I L R L M M �Q �Q R R L U �U V V X X V X Y Y �[ �[ \ \ �^ �^ _ _ �a a b b �d d e e �g g h h �j j k k �m m n n �p 	p q q �t t u u v v w w x x y y z �z { �{ | | !} } *~ ~ ,  /� � 3� � 8� � >� � E� t� � W� � -� � ,� � � �� � �� � M� � U� � \� � b� � g� � k� � n� � p� �� � +� � � � � }� � � � � z� � � � �   � � � � �   � � � � �   � � � � �   � � � � � � �� � �� � �� �   � � �� �   � � �� �   � v� � � � � �� � � � � � � � � y� � |� � ~� � u� � � � � �� � � � � � � �� � �� � �� � �� � �� � �� � �� � � �� �   � � �� � � � � �� �� � � ��  � � � �� � � � �� � � �  � � � � � � � � � �� �  � � �� � �� ��� 2 � � � � � � � E� 	� IJ� G 5 C� �Dg�j� #',($!qwrx"""0s{&&&/&89+� &� .� .).%1171:1>1AB-626*"X939Y9|ut=4=Z^{@5[XC1BD FF
HDHFK� 1 ��v�F N}MOhOkOnOqOtO~Ow\y6� X;X?@W@\[O^_=]_i_l_o_r_u__x]/ gPg`�jQja�mRmb��pSpc��sTsd��vVvfL�O0 {� {<=z}U}eN�� �K4 H3 � � � �B ��g�& �A ��j�' �@ m�p�m�p�( ��? ) �G �s�s�}�* �v�+ �E L, �I ����Y �M �\ �_ �b �q �n �k �h �e �U ����Q ���������� ���������������������������� ����������������������������
��� ��[ ���������������{ ��������������������������� ������^ ��������������z �a 	�������y p ������x 
m �����w j g ����v ��u �d �t ���� | ""+"-"0"4"9"?"FM!*#} N,$,O~ V/%/P/W ]3&3Q3X3^� c8'8R8Y8_8d� h>(>S>Z>`>e>i� lE)ETE[EaEfEjEm� o� "N.N1N5N:N@NGU*� NV2V6V;VAVH\,� V]7]<]B]Ib/� ]c=cCcJg3� chDhKk8� hlLn>� lpE� oy|.~69z� &w� vz� qx� }"� r{� � s������ ����� ���� ��� � ���� ��� ����� � ������  ���� ���� �� �� � ��� ���� �� �� �� �� ��� � �  D          �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 