��  CCircuit��  CSerializeHack           ��  CPart          ���  CLED_G�� 	 CTerminal  p�q                �          
�  pq1                            d�         ��      ��  COR
�  Hh]i               �          
�  Hx]y               �          
�  tp�q               �            \dt|           ��    �� 	 CResistor��  CValue  ����    330          �t@      �?   
�  ����                �          
�  ����               �            ����         ��      ��  CAND
�  `�u�               �          
�  `�u�              @          
�  ����               �            t���           ��    �
�  ���               �          
�  ���     	          �          
�  $�9�               �            �$�           ��    �� 	 CInverter
�  �               �          
�  $9              @            $     #      ��    ��  ���    300          �r@      �?   
�  ��                �          
�  �     
          �            ��     '    ��      ��  c���    330          �t@      �?   
�  ����      	          �          
�  ���               �            ����     +    ��      ��  CEarth
�  ����                             ����     /    ��      ��  CBattery�  #IKW    5V(          @      �? V 
�  X0YE               @          
�  X\Yq                            LDd\     3    ��      -�
�  X�Y�                             K�c�     6    ��      ��  ����    330          �t@      �?   
�  ����                �          
�  ���	               �            ����     9    ��      ��  CLED
�  (=      
          �          
�  Ti                            <,T     =    ��      ��  CLED_Y
�  �(�=                �          
�  �T�i                            |<�T     A    ��      �
�  �(�=                �          
�  �T�i                            �<T     D    ��      ��  CSPST��  CToggle  H8h      G   
�  dy               �          
�  8M               @            Ld    J      ��    F�H�  �H�h      L   
�  �d�y     	          �          
�  �8�M               @            |L�d    N      ��    F�H�  �Hh      P   
�  �d�y               �          
�  �8�M               @            �L�d    R      ��              ���  CWire  ����       U�  �h��       U�  ��I�      U�  H�I1       U�  H0q1      U�  p�q�       U�  p���      U�  �xIy      U�  �hi      U�  �p��       U�  �p�q      U�   hIi      U�   8!i       U�   8�9      U�  ���9       U�  ���y       U��� 
 CCrossOver  ��      g�  ~���        ����      U�  ����       U�g�  ��        ��       U�g�  ~���        ����      	 U�  ����       U�  ��)       U�  ����       U�  `�a       U�  8a      U�  `�a�       U�  8�a�      U�  ��      U�  ���       U�  ���      U�g�  |�      g�  ��        x�       U�  ����      	 U�  ����      	 U�  ����     	 U�g�  ��        ����     	 U�g�  ~|��        �x��      	 U�g�  |�      g�  ~|��        ����      U�  �x��       U�  ()     
 U�   )      
 U�  � �)       U�  ����     	 U�  ����      U�  �h�i      U�  XpY�       U�  �0�9       U�  X0�1      U�  �8�9      U�  �89                �                     [    Z  a   ]    `  _    \  t   r    d  q   }      u # v # $ $ s ' k ' ( ( � + � + , , � / � / 3 � 3 4 4 � 6 � 6 9 o 9 : : p = � = > > ^ A � A B B � D p D E E W J J y K � K N N � O � O R R � S � S W � � X V Y X Z Y  \  [  e  B > `   _ b  c a b d  c f ] f l f n o e � f k h y ' m i � � j 9 : D �   s $ r u    t w # x v k w y � y � J x  ~  ~ | }  { m | � � N  � z � � j q R � � = ( � , A m + / V E ^ 4 6 � S 3 � � O � K             �$s�        @     +        @            @    "V  (      �8                
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 