��  CCircuit��  CSerializeHack           ��  CPart    0   0     ���  CAND�� 	 CTerminal  lP�Q              @          
�  l@�A               �          
�  @HUI               �            T<lT          ��    ��  CEarth
�  � �       	          W�/�1�?    ��         ��      ��  CClock
�  D � Y �               @            , � D �          ����     �� 	 CVoltRail��  CValue  + q S      5V(          @      �? V 
�  \ x q y               @            T t \ |          ����     ��  CSPST��  CToggle  � � � �         
�  p x � y       	       @          
�  � x � y               @            � t � |           ��    �� 
 CCounter10
�  x -y               @          
�  � -�               @          
�  @� A�                �          
�  L� a�                �          
�  L� a�               @          
�  L� a�                �          
�  Lp aq                �            ,l L�      !      ��  ,   �� 	 CPushMake��  CKey  J� n�       )   
�  @� A�               @          
�  @� A�        	        �            8� D�     ,      ��    ��  C4511
�  �p �q                �          
�  �� ��                �          
�  �� ��               @          
�  �� ��                �          
�  �� ��               @          
�  �� ��               @          
�  �� ��               @          
�  �� ��                �          
�  �� ��                �          
�  �� ��         {��.@�W�/�1��  
�  �� ��         {��.@�W�/�1��  
�  �� ��                �          
�  �� ��         {��.@�W�/�1��  
�  �p �q      
   {��.@�W�/�1��    �l ��      0      ��  h   �� 
 CResistors�  �^ l     220        �k@      �?   
�  �p �q      
 	 {��.@�W�/�1�?  
�  �� ��       	 {��.@�W�/�1�?  
�  �� ��       	        �          
�  �� ��       	 {��.@�W�/�1�?  
�  �� ��       	 {��.@�W�/�1�?  
�  �� ��       	        �          
�  �� ��       	        �          
�  �� ��                �          
�  � !�                �          
�  � !�                �          
�  � !�                �          
�  � !�         �i�n� @�W�/�1��  
�  � !�         �i�n� @�W�/�1��  
�  � !�      	          �          
�  � !�         �i�n� @�W�/�1��  
�  p !q         �i�n� @�W�/�1��    �l �      A      �� v   ��  CSevenSegmentDisplay
�  p� ��         �i�n� @ W�/�1�?  
�  p� ��         �i�n� @ W�/�1�?  
�  p� ��                �          
�  p� ��                �          
�  �� �                 W�/�1��  
�  �� ��                �          
�  �� ��         �i�n� @ W�/�1�?  
�  �� ��         �i�n� @ W�/�1�?  
�  �� ��      	          �            �� ��      S 	     ��0 <                0   0     ���  CWire  �PQ      ]�   H Q       ]�  �H I       ]�  �P �Q       ]��� 
 CCrossOver  ~l �t       c�  ~| ��         �H ��        ]�  `� ��       ]�  �P �q        ]�c�  ~l �t         `p �q       ]�c�  ~| ��         `� ��       ]�  �� ��       ]�  �@�A      ]�  �P �A       ]�  �p �q       ]�  0� A�       ]�c�  .� 4�       c�  .4      c�  .4        0� 1I       ]�  0HAI      ]�c�  .� 4�          � A�       ]�c�  .4        � y	      ]�c�  .4        � �      ]�   � Y�       ]�   � a�       ]�  � x � y       ]�c�  � � �       c�  � � � �         � � �       ]�  � �        ]�c�  � � �       c�  � � �          x �        ]�c�  � � � �       c�  � � � �         � x � 	       ]�  � � � �        ]�  X � � �       ]�  � � �        ]�  � x y       ]�   x y       ]�  `� ��       ]�   � ��      	 ]�  �� ��       	 ]�  �� ��       ]�   � ��       ]�  �� ��        ]�   p �q       ]�  �p ��        ]�  �� ��       ]�   � q�       ]�  p� q�        ]�   � i�       ]�  h� i�        ]�  h� q�       ]�  `� a�        ]�  `� q�       ]�  X� q�       ]�  X� Y�        ]�  x� y	       ]�  x� ��       ]�  x� y�        ]�  x� ��       ]�  �� ��       ]�  �� �       ]�c�  � � � �       c�  � � �         � � �           0   0     �    0   0         0   0       ^   m  u   W    �         ~ ! � ! " � " # # - $ $ � % % f & & j ' ' h , , v - p - 0 o 0 1 j 1 2 l 2 3 � 3 4 � 4 5 � 5 6 � 6 7 7 G 8 8 F 9 9 E : : D ; ; C < < B = = A A = A B < B C ; C D : D E 9 E F 8 F G 7 G H   H I I   J J | K K } L L � M M � N N � O O � P P � S � S T � T U � U V � V W W  X X   Y Y � Z Z � [ [ �  _ ` ^ b _ g n b i b k ` l % b a o h d ' g j e & 1 f 2  n a m h 0 q # q w q y q { p u q  v r � , x s � � z t � � J � K �  �  �  � � "  � � � � � � v � � � � ~ x  �  � � z � � � ! $ 3 N � � [ Z � O � � � P � � � Y � M � � S L � � � � T } � � U � V | � � x � 4 � � � 5 � 6 � z � � � � � �            �$s�        @     +        @            @    "V  (      �P                
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 