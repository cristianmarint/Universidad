��  CCircuit��  CSerializeHack           ��  CPart              ��� 	 CInverter�� 	 CTerminal  Pe     
          �          
�  |�              @            d|           ��    ��  COR
�  � �               �          
�  ��              @          
�  )	        ���P�p@����\*��    ��            ��    ��  CAND
�  �� ��               @          
�  �� ��                �          
�  �� ��                �            �� ��            ��    �
�  `� u�               @          
�  `� u�               @          
�  �� ��               @            t� ��            ��    �
�  � �                �          
�  4� I�               @            � 4�            ��    �
�  �� ��                �          
�  � !�               @            �� �            ��    �� 	 CResistor��  CValue  K�k�    330          �t@      �?   
�  ppq�         ���P�p@����\*�?  
�  p�q�        �٭$M� @����\*��    l�t�     %    ��      ��  CLED_G
�  pq         �٭$M� @����\*�?  
�  p4qI                ����\*��    d�4     )   ��      ��  CSPST��  CToggle  Xx x�       ,   
�  P� Q�      
          �          
�  Ph Q}                @            L| T�     /      ��    +�-�  �x ��       1   
�  �� ��                �          
�  �h �}                @            �| ��     3      ��    +�-�  �x �       5   
�  �� ��                �          
�  �h �}                @            �| ��     7      ��    +�-�  p 0�       9   
�  � 	�                �          
�  ` 	u                @            t �     ;      ��    ��  CBattery#�   � 3 �     5V(          @      �? V 
�  @ � A �                @          
�  @ A                             4 � L      @    ��      ��  CLED_Y
�  PQ                �          
�  P4QI                            Dd4     D    ��      B�
�  ��      	          �          
�  �4�I                            ��4     G    ��      B�
�  � �                �          
�  �,�A                            ��,     J    ��      B�
�   	                �          
�  ,	A                            � ,     M    ��      !�#�  +�K�    330          �t@      �?   
�  PxQ�      
          �          
�  P�Q�               �            L�T�     Q    ��      !�#�  ����    330          �t@      �?   
�  �x��                �          
�  ����     	          �            ����     U    ��      !�#�  ����    330          �t@      �?   
�  �x��                �          
�  ����               �            ����     Y    ��      !�#�  � ��    330          �t@      �?   
�  x	�                �          
�  �	�               �            ��     ]    ��      ��  CEarth
�  @ �A �                 ����\*�?    3 �K �     a    ��                    ���  CWire  pqq       c�  (q	      c�  �� ��       c�  �� �       c�  ��      c��� 
 CCrossOver  N� T�       j�  N� T�       j�  N� T�         P� Q      
 c�  PQy      
 c�  � �i        c�  �� ��        c�j�  N� T�         �� ��       c�j�  �� ��       j�  �� ��         �� ��        c�  �� �y       c�  �� ��        c�  `� a�        c�j�  N� T�       j�  �� ��          � a�       c�  `� a�        c�j�  N� T�       j�  �� ��       j�  �� ��         H� a�       c�  � 	�        c�  � 	y       c�j�  �� ��         �� ��        c�  �� �y       c�   	a        c�  PHQ�       c�  P�q�      c�  pHq�       c�  p�q	       c�   �       c�  P Qi        c�  � Q       c�  � �i        c�  � �       c�  @  	       c�  @  A �        c�  X �q �      c�  @ �Y �      c�  X �Y �       c�  @ �Y �      c�  @ A �       c�  @ �A �       c�  ����      c�  ��Q�      c�  ���      c�  �H��       c�  @	�       c�  �@��       c�  p �q �       c�  p �	�      c�  P�Q	       c�  ���	      	 c�  ���       c�  �	                     �                             n    h  g   h    e  w   p    f  |   x    w  �    }  �      y % d % & & � ) � ) * * � / / i 0 � 0 3 3 s 4 � 4 7 7 � 8 o 8 ; ; � < � < @ � @ A A � D � D E E � G � G H H � J � J K K � M � M N N � Q n Q R R � U v U V V � Y � Y Z Z � ] � ] ^ ^ � a � a e %  d  g f    i ~ i z i r /  i Q � 8  q q m v p s  s { 3 q s U    y y l y u   x  } } k } t } �  | ;  � ] � � 7  � Y � < E � � � * � & ) � � � 0 � � � 4 o � � � � @ � � � � � � � � A � � a � � � � � � H � N � K � � � � � R D V G Z J ^ M             �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 