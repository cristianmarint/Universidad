��  CCircuit��  CSerializeHack           ��  CPart    0   0     ���  CEarth�� 	 CTerminal  � �       	          W�/�1�?    ��         ��      ��  CClock
�  D � Y �                             , � D �          ����     �� 	 CVoltRail��  CValue  + q S      5V(          @      �? V 
�  \ x q y               @            T t \ |          ����     ��  CSPST��  CToggle  � � � �         
�  p x � y       	       @          
�  � x � y               @            � t � |           ��    �� 
 CCounter10
�  x -y               @          
�  � -�                           
�  @� A�                �          
�  L� a�                �          
�  L� a�                �          
�  L� a�                �          
�  Lp aq               @            ,l L�            ��  ,   �� 	 CPushMake��  CKey  J� n�       $   
�  @� A�               @          
�  @� A�        	        �            8� D�     '      ��    ��  C4511
�  �p �q               @          
�  �� ��                �          
�  �� ��                �          
�  �� ��                �          
�  �� ��               @          
�  �� ��               @          
�  �� ��                           
�  �� ��                �          
�  �� ��                �          
�  �� ��                �          
�  �� ��                �          
�  �� ��                �          
�  �� ��         {��.@�W�/�1��  
�  �p �q      
   {��.@�W�/�1��    �l ��      +      ��  h   �� 
 CResistors�  �^ l     220        �k@      �?   
�  �p �q      
 	 {��.@�W�/�1�?  
�  �� ��       	 {��.@�W�/�1�?  
�  �� ��       	        �          
�  �� ��       	        �          
�  �� ��       	        �          
�  �� ��       	        �          
�  �� ��       	        �          
�  �� ��                �          
�  � !�                �          
�  � !�                �          
�  � !�                �          
�  � !�                �          
�  � !�                �          
�  � !�      	          �          
�  � !�         �i�n� @�W�/�1��  
�  p !q         �i�n� @�W�/�1��    �l �      <      �� v   ��  CSevenSegmentDisplay
�  p� ��                �          
�  p� ��                �          
�  p� ��                �          
�  p� ��                �          
�  �� �                 W�/�1��  
�  �� ��                �          
�  �� ��         �i�n� @ W�/�1�?  
�  �� ��         �i�n� @ W�/�1�?  
�  �� ��      	          �            �� ��      N 	     ��0 <                 0   0     ���  CWire  � �      X��� 
 CCrossOver  � � �       [�  � � � �         � � �       X�  � �        X�[�  � � �       [�  � � �          x �        X�[�  � � � �       [�  � � � �         � x � 	       X�  � � � �        X�  X � � �       X�  � � �        X�  � x y       X�  � x � y       X�   x y       X�   � A�       X�  `p �q       X�  `� ��       X�  `� ��       X�  `� ��       X�   � ��      	 X�  �� ��       	 X�  �� ��       X�   � ��       X�  �� ��        X�   p �q       X�  �p ��        X�  �� ��       X�   � q�       X�  p� q�        X�   � i�       X�  h� i�        X�  h� q�       X�   � a�       X�  `� a�        X�  `� q�       X�  X� q�       X�  X� Y�        X�   � Y�       X�  � y	      X�  x� y	       X�  x� ��       X�  x� y�        X�  x� ��       X�  �� ��       X�  �� �       X�[�  � � � �       [�  � � �         � � �           0   0     �    0   0         0   0      R    f         i  j   ^    (   o     n ! ! m " " l ' ' k (  ( + l + , m , - n - . o . / � / 0 � 0 1 � 1 2 2 B 3 3 A 4 4 @ 5 5 ? 6 6 > 7 7 = 8 8 < < 8 < = 7 = > 6 > ? 5 ? @ 4 @ A 3 A B 2 B C   C D D   E E � F F } G G z H H x I I p J J s K K u N y N O | O P  P Q � Q R R  S S   T T w U U r V V q g � Z ` Z c e  Z � _ \ _ � j k b ] b � i � Z f  e � Y b _  h h  _ ' " + ! ,   -  . I q p V U t J t s r K v u w T v H y x N G { z | { O F ~ }  ~ P � Q � � E � b � � � � / � � � 0 � 1 � Y � d � a g ^            �$s�        @     +        @            @    "V  (      �P                
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 