��  CCircuit��  CSerializeHack           ��  CPart    0   0     ���  CECapacitor��  CValue  � ��    100�F(    -C��6?      �?�F �� 	 CTerminal   p!�      !   �H���?ʒ)d,`�  �   �!�     "           ʒ)d,`?    �,�        ��      q��gC��>��  CLED_G�  � �!               �          �  � �!     "                       ��4        ��      ��  �@�A               �          �  �@�A     "                       �4�T        ��      ��  �`�a               �          �  �`�a     "                       �T�t        ��      ��  ����               �          �  ����     "                       �t��        ��      ��  ����                �          �  ����     "                       ����        ��      ��  � �               �          �  � �     "                       �� �         ��      ��  �� ��                �          �  �� ��      "                       �� ��     #    ��      ��  �� ��                �          �  �� ��      "                       �� ��     &    ��      ��  �� ��         B��� @ �:�?  �  �� ��      "            �:��    �� ��     )  
 ��      ��  �� ��                �          �  �� ��      "                       �t ��     ,    ��      �� 
 CResistors
�  0P$    220        �k@      �?   �   (5)               �          �   859               �          �   H5I               �          �   X5Y     
          �          �   h5i               �          �   x5y               �          �   �5�               �          �   �5�               �          �  L�a�               �          �  L�a�               �          �  Lxay               �          �  Lhai               �          �  LXaY               �          �  LHaI     	          �          �  L8a9                �          �  L(a)               �            4$L�     1      �� v   .�
�  0n P|     220        �k@      �?   �   � 5�       	        �          �   � 5�       	 �v��D/@'�:�?  �   � 5�       	        �          �   � 5�       	        �          �   � 5�       	        �          �   � 5�       	        �          �   � 5�       	        �          �   � 5�       	        �          �  L� a�                �          �  L� a�                �          �  L� a�                �          �  L� a�                �          �  L� a�                �          �  L� a�                �          �  L� a�         B��� @'�:��  �  L� a�                �            4| L�      C      �� v   ��  CDecoder�  �� ��      ) 	       @          �  �� ��      ( 	        �          �  �� ��      ' 	        �          �  �� ��      & 	        �          �  �� �	               �          �   � 	               �          �  � !�                �          �  � !�                �          �  � !�                �          �  � !�                �          �  � !�                �          �  � !�                �          �  � !�         �v��D/@@�:��  �  � !�                �            �| �      U      ��  T   �� 	 CResistor
�  � � �     470          `}@      �?   �   � !�       #         @<s���?�?  �   � !	     -   �H���?<s���?��    � $�      f    ��      �� 
 CVResistor��  CSlider  0?<     
�  � !/    0k     F]t�1�@        k 
   l �   !      - 	 �H���?Ȓ)d,`�  �   4!I     !   �H���?Ȓ)d,`?    ,4     m    ��      ��  C555�  �� ��       #         @N贁Nk?  �  �� ��       #         @          �  �� ��      -   �H���?��8��J�?  �  �� ��      !   �H���?          �  � �     !   �H���?          �  ��     "           ao9 ?��  �  ��     .   ������
@       �  �  �� 	�      $          �            �� �     q    ��   (   ��  CEarth�   �!�      "           �Hi�Ϗ�?    �+�     {    ��      ��    !5      $          �          �   L!a     ,          �            44L     }    ��      c�
�  �y�    220          �k@      �?   �   `!u      , 	        �          �   �!�     "                       t$�     �    ��      ��  CSPST��  CToggle  � � � �      �   �  � � � �      *         @z(=e�?  �  � � � �      #         @z(=e��    � � � �      �     ��    y��  P � Q �       + 	         z(=e��    C � [      �    ��      ��  CBattery
�   � C �     5V(          @      �? V �  P � Q �       *         @z(=e��  �  P � Q �      +           z(=e�?    D � \ �      �    ��      �� 	 CPushMake��  CKey  �� �      �   �  ��)     #         @          �  �� ��       % 	        �            �� �    �      ��    �� 
 CCounter10�  �� ��      #         @          �  �� ��      $          �          �  �� ��      %          �          �  �� ��      &          �          �  �� ��      '          �          �  �� ��      (          �          �  �� ��      )         @            �� ��      �      ��  ,       0   0     ���  CWire   �!�      " ��   ���     " ��  ����      " ��  ����      " ��  �`��      " ��  �@�a      " ��  � �A      " ��  � �!      " ��  �� �      " ��  �� ��       " ��  �� ��       " ��  �� ��       " ��  � �!      ��  �� �!       ��  `� ��       ��  �� �       ��  �� ��        ��  �� �A       ��  � �      ��  `� ��       ��  �� ��       ��  h���       ��  h8i�        ��  `8i9       ��  p���      ��  p(q�       ��  `(q)      ��  x`�a      ��  x� ya       ��  `� y�       ��  �@�A      ��  `� ��       ��  `� ��       ��  �� ��        ��  �� ��       ��  `� ��       ��  �� ��        ��  `� ��       ��  `� ��       ��  �8!9      ��  ��9       ��   (!)      ��   )       ��   � ��      # ��  � !�      $ ��   � !�       # ��  �� ��       # ��  �� ��      # ��  �� ��       # ��  p� ��      - ��  p� q	      - ��  �� ��      ! ��   `�a     ! ��   H!a      ! ��   `!q      ! ��   q	     - ��  � �     ! ��  �� �      ! ��  � �a      ! ��   � !!      $ ��   �!�      " ��   �!�      " ��  P � � �      * ��  � � !�      # ��  ���      " ��   ���     " ��  x(�)     # ��  �� y�      # ��  ��!�     " ��  x� ��      # ���� 
 CCrossOver  v� |�         x� y)      # ���  v� |�          � ��      $ ��  �� ��       $     0   0     �    0   0         0   0      �    �  �    �  �    �  �    �  �    �  �    �   �   ! ! � # � # $ $ � & � & ' ' � ) � ) * * � , � , - - � 1 � 1 2 � 2 3   3 4   4 5   5 6   6 7   7 8   8 9 9   : :   ; ;   < <   = =   > >   ? ? � @ @ � C b C D a D E ` E F _ F G ^ G H ] H I \ I J [ J K K � L L � M M � N N � O O � P P � Q Q � R R � U � U V � V W � W X � X Y Y � Z Z � [ [ J \ \ I ] ] H ^ ^ G _ _ F ` ` E a a D b b C f � f g g � m g m n n � q � q r � r s � s t � t u � u v v � w w   x x � { � { } � } ~ ~ � � ~ � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � X � � W � � V � � U � � � �  �  �  �  �  � ! � $ � ' � * � - � �  � � M � � � � � � � �   N � � # �  � � ? � �  � � @ � �  � � K � �  L � O � � � � & P � � ) Q � R , � 2 Y � � 1 Z � � � x � � f � r � � � q � s � � � t � � n � �  m � � u � � � � � }  � � { � � � � v � � � � � � � � � � � � � � � � � � � � �  /          �$s�        @     +        @            @    "V  (      �P                
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 