��  CCircuit��  CSerializeHack           ��  CPart�� 
 CTextLabel  1�Y�    Decodi.      �  �� �     CI 555 generador de pulsos          0   0     ���  CECapacitor��  CValue  ���    100�F(    -C��6?      �?�F �� 	 CTerminal  ��         �[F2���?t�6�o�9�  �  �     
           t�6�o�9?    ��        ��      �O4]�"?�� 	 CPushMake��  CKey  H� l�          �  8� M�      $         @          �  d� y�                �            L� d�            ��    ��  CAND�    5                �          �  � �5               @          �  �L�a               �            �4L          ��    �� 
 CResistors�  1�Q�    220          �k@      �?   �  ����      " 	 |��.@�W�/�1�?  �  ����      4 	 {��.@�W�/�1�?  �  ����       	 |��.@�W�/�1�?  �  ����       	        �          �  ����       	 |��.@�W�/�1�?  �  x�y�       	 |��.@�W�/�1�?  �  h�i�      . 	 |��.@�W�/�1�?  �  X�Y�                �          �  X�Y               �          �  h�i     9   �i�n� @�W�/�1��  �  x�y     8   �i�n� @�W�/�1��  �  ���     7   �i�n� @�W�/�1��  �  ���     6          �          �  ���     !   �i�n� @�W�/�1��  �  ���        �i�n� @�W�/�1��  �  ���     ;   �i�n� @�W�/�1��    R���           �� v   ��  CSevenSegmentDisplay�  p@�A     6          �          �  pP�Q     7   �i�n� @ W�/�1�?  �  p`�a     8   �i�n� @ W�/�1�?  �  pp�q     9   �i�n� @ W�/�1�?  �  �|��     5           @A�c=岿  �  �p�q     :          �          �  �`�a     ;   �i�n� @ W�/�1�?  �  �P�Q        �i�n� @ W�/�1�?  �  �@�A     !   �i�n� @ W�/�1�?    �<�|     2 	     ��0 <           ��  CEarth�  ����      5 	         @A�c=�?    ����     =    ��      ;��  � �                              � $�     ?    ��      ;��  H�I�      3 	         @A�c=�?    ;�S�     A    ��      0��   H5I     /          �          �   X5Y               �          �   h5i               �          �   x5y     %          �          �  H�I�     3           @A�c=墿  �  dxyy     &          �          �  dhyi     2   �i�n� @ W�/�1�?  �  dXyY     1   �i�n� @ W�/�1�?  �  dHyI     0   �i�n� @ W�/�1�?    4Dd�     C 	     ��0 <             ��  ���    220          �k@      �?   �  x�y�      ' 	 |��.@�W�/�1�?  �  h�i�      ( 	 |��.@�W�/�1�?  �  X�Y�      ) 	 |��.@�W�/�1�?  �  H�I�      * 	        �          �  8�9�      + 	        �          �  (�)�      , 	        �          �  ��      - 	        �          �  �	�                �          �  �		               �          �  �	     %          �          �  (�)	               �          �  8�9	               �          �  H�I	     /          �          �  X�Y	     0   �i�n� @�W�/�1��  �  h�i	     1   �i�n� @�W�/�1��  �  x�y	     2   �i�n� @�W�/�1��    �|�    N      �� v   ��  C4511�  x�y�               @          �  h�i�               @          �  X�Y�               @          �  H�I�                �          �  8�9�      $         @          �  (�)�      $         @          �  ��                            �  ��     -          �          �  (�)�     ,          �          �  8�9�     +          �          �  H�I�     *          �          �  X�Y�     )   |��.@�W�/�1��  �  h�i�     (   |��.@�W�/�1��  �  x�y�     '   |��.@�W�/�1��    �|�    `      ��  h   ^��  �x��                �          �  �x��                �          �  �x��                �          �  �x��                �          �  �x��      $         @          �  xxy�      $         @          �  hxi�                            �  h�i�     .   |��.@�W�/�1��  �  x�y�        |��.@�W�/�1��  �  ����        |��.@�W�/�1��  �  ����               �          �  ����        |��.@�W�/�1��  �  ����     4   {��.@�W�/�1��  �  ����     "   |��.@�W�/�1��    `���    o      ��  h   �� 
 CCounter10�  ��-      $         @          �  ��-                �          �  �@�A               �          �  �L�a               �          �  �L�a               �          �  �L�a               �          �  �L�a               �            �,�L          ��  ,   }��  pq-      $         @          �  PQ-                �          �  0@EA               �          �  HLIa               �          �  XLYa              @          �  hLia              @          �  xLya              @            D,|L    �      ��  ,   ��  CBattery�  !3/    5V(          @      �? V �  @A               @���Z�$��  �  @4AI                ���Z�$�?    4L4     �    ��      ;��  @HA]       	         ���Z�$��    3\Kd     �    ��      ��  CSPST��  CToggle  ��0     �   �  ��	              @���Z�$�?  �  ��	     $         @���Z�$��    ��     �     ��    �� 	 CResistor�  ���    220          �k@      �?   �  ��       	        �          �  �     
                       ��     �    ��      ��  CLED_G�  ��                �          �  ��               �            �$�     �    ��      ;��  �x��       	         ?�����?    ����     �    ��      ;��  (=      
           t�6�o�9�    <D     �    ��      ��  C555�  �(�=      $         @N贁Nk?  �  �(�=      $         @          �  �@�A     	   ������?l��k-�?  �  �P�Q        �[F2���?          �  �`�a        �[F2���?          �  �d�y                ?�����  �  �d�y        ������
@       �  �  �P�Q               �            �<�d     �    ��   (   �� 
 CVResistor��  CSlider   t/�     �  ���    3.33k     �����F�@�������?k 
   � �  h}      	 	 ������?u�6�o�9�  �  ��        �[F2���?u�6�o�9?    |�     �    ��      ���  �AO    470          `}@      �?   �  (=      $         @��]�	Q�?  �  Ti     	   ������?��]�	Q��    <T     �    ��          0   0     ���  CWire�� 
 CCrossOver  ~�      ��  ~�        �� �A       ��  x� ��       ����  ~�      ��  .4      ��  ��      ��  ��      ��  6<      ��  v|      ��        ��  ��        Q      ����  ~�      ��  ��        x�	     $ ����  � �         �� 1�       ����  .4      ��  .4      ��  .4        0� 1A       ����  .4      ��          �9      ����  .4      ��  ��      ��  6<      ��          �q	     $ ��  8 �      ����  � �       ��        ��  $      ��        ��          � i        ��   � 9�      $ ��   � !	      $ ��  �!	     $ ��   y	     $ ����  ��      ��  ��        �� �       ��  �� ��       ����  ��      ��  ��        �� �a       ��  �`�a      ����  vl|t        xhy�       ��  x`yi       ����  �d�l        xh�i      ����  �d�l        ��q      $ ��  � �i       ����  6<      ��  6<        8 9       ��  ��!       ����  $          !!      ��   `Ia      ��    !a       ����  �d�l        �`�y      $ ����  �d�l      ��  �d�l      ��  �d�l      ��  �d�l      ��  �d�l        hhi       ��  x`�a     $ ����  v|        xya      $ ��  xx�y     $ ��  h�        ��  hhiy        ����  �d�l        �`�y       ����  �d�l        �`�y       ����  �d�l        �`�y       ����  �d�l        �`�y       ��  �`�a     ; ��  � �     ; ��  � �       ��  ��      ��  � �a      ; ��  �P�Q      ��  � �      ! ��  ��     ! ��  ��Q       ��  ��A      ! ��  �@�A     ! ��  � �1      6 ��  h0�1     6 ��  h0iA      6 ��  h@qA     6 ��  `PqQ     7 ��  `(aQ      7 ��  � �)      7 ��  X`qa     8 ��  X Ya      8 ��  `(�)     7 ��  X y!     8 ��  x y!      8 ��  Ppqq     9 ��  PQq      9 ��  Pi     9 ��  h i      9 ��    y      % ��  p`�a      ��  (�9�     $ ��  8p9�      $ ��  p�	     $ ��  pq      $ ����  vl|t      ��  fllt      ��  Vl\t      ��  FlLt        8p�q     $ ����  fllt        h`i�       ����  Vl\t        X`Y�       ����  FlLt        H`I�       ��  !      % ��    !     % ��   x!y     % ��  ())       ��  ())      ��  091      ��  (	i       ��  h!i      ��  891       ��  0Y       ��  X!Y      ��  H!I     / ��  8I      / ��  8I9     / ��  HI9      / ��  xH�I     0 ��  � �I      0 ��  ��Y      1 ��  X �!     0 ��  XY!      0 ��  xX�Y     1 ��  ��i      2 ��  h�     1 ��  hi      1 ��  x�	     2 ��  xh�i     2 ��  @�	      ��  �	     $ ��  PQ       ��  Q       ����  ��        ��      $ ��  �	     $ ��  )      
 ��        
 ��       
 ��         
 ��  P�       ��  �PQ      ��  p`q�       ��  pPqa       ��  hai     	 ��  ��       ��  ��       ��  �q�      ��  pP�Q      ��  `@ai      	 ��  `@�A     	 ��  ��)      $ ��  ��	     $ ��  ��)      $ ��  )      $     0   0     �    0   0         0   0      m   e �    �  �   �    �   |   ! { ! " z " # y # $ x $ % w % & v & '   ' ( (   ) ) 1* * -+ + (, , "- - . . / / 2 %2 3 &3 4 )4 5 .5 6 6 = 7 7   8 8 9 9 : : != 6 = ? ? � A G A C NC D MD E JE F EF G G A H H   I I \J J WK K RN m N O l O P k P Q j Q R i R S h S T g T U   U V V   W W CX X FY Y KZ Z Q[ [ V\ \ Z] ] [` � ` a =a b ?b c Ac d 5d e 4e f f g g T h h S i i R j j Q k k P l l O m m N o o p p q q r r s s t t u u v v & w w % x x $ y y # z z " { { ! | |    a � � � � � � � � � � � � � � � 7� � _� � � � � � A� � ?� � =� � � � ]� � � � � � � � ]� � � ^� � � � � g� h� � � � � � � � d� � s� � u� � r� � p� � 3� � � � � �   � � i� � � � � n� v� � � l� � � � � �  � � � � � � � � � � � � � � � b`_� � � � � a� � � � � � � � � � � � � � � � � � � � � � � � � � � 7� � � � � � � � � � � � ? �  � � s� � 
� � � � � � � � � � � � � � �  � 9� ` � � � � � � � � 68� � � � � � � � �  � �    � � � 	s 

� � 	t � f u � o � p � q � r 8 / . 9 -  !:  , #$"#%$2 '3 +&+ +*4 ,)'(*-* ,/5 0./1) 0DEj� e d 84� � 6� 8� 8>8@8B5� =:� a ?;� b A<� c W D2C2F X GIFLKGJIE Y HHMLD OC PNOQZ PK SURYWVS[ UJ T[\ZT\ Y] XI X� � � c� � � ia� �  vte�  fdg� f`� � hkop3� qn � omjk� rlq� t� u� c� ^�  <          �$s�        @     +        @            @    "V  (      �P                
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 